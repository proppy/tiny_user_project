magic
tech sky130A
magscale 1 2
timestamp 1662467768
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 1104 2128 49666 47376
<< metal2 >>
rect 662 49200 718 50000
rect 12898 49200 12954 50000
rect 25134 49200 25190 50000
rect 37370 49200 37426 50000
rect 49606 49200 49662 50000
rect 18 0 74 800
rect 12254 0 12310 800
rect 24490 0 24546 800
rect 36726 0 36782 800
rect 48962 0 49018 800
<< obsm2 >>
rect 1398 49144 12842 49314
rect 13010 49144 25078 49314
rect 25246 49144 37314 49314
rect 37482 49144 49550 49314
rect 1398 856 49660 49144
rect 1398 800 12198 856
rect 12366 800 24434 856
rect 24602 800 36670 856
rect 36838 800 48906 856
rect 49074 800 49660 856
<< metal3 >>
rect 0 38088 800 38208
rect 49200 37408 50000 37528
rect 0 25168 800 25288
rect 49200 24488 50000 24608
rect 0 12248 800 12368
rect 49200 11568 50000 11688
<< obsm3 >>
rect 800 38288 49200 47361
rect 880 38008 49200 38288
rect 800 37608 49200 38008
rect 800 37328 49120 37608
rect 800 25368 49200 37328
rect 880 25088 49200 25368
rect 800 24688 49200 25088
rect 800 24408 49120 24688
rect 800 12448 49200 24408
rect 880 12168 49200 12448
rect 800 11768 49200 12168
rect 800 11488 49120 11768
rect 800 2143 49200 11488
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< labels >>
rlabel metal3 s 49200 24488 50000 24608 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 662 49200 718 50000 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 49200 37408 50000 37528 6 io_in[2]
port 3 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 io_in[3]
port 4 nsew signal input
rlabel metal2 s 25134 49200 25190 50000 6 io_in[4]
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_in[5]
port 6 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 io_in[6]
port 7 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 io_in[7]
port 8 nsew signal input
rlabel metal2 s 37370 49200 37426 50000 6 io_out[0]
port 9 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_out[1]
port 10 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 io_out[2]
port 11 nsew signal output
rlabel metal2 s 49606 49200 49662 50000 6 io_out[3]
port 12 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_out[4]
port 13 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_out[5]
port 14 nsew signal output
rlabel metal2 s 12898 49200 12954 50000 6 io_out[6]
port 15 nsew signal output
rlabel metal3 s 49200 11568 50000 11688 6 io_out[7]
port 16 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 596062
string GDS_FILE /home/runner/work/tiny_user_project/tiny_user_project/openlane/user_module/runs/22_09_06_12_34/results/signoff/user_module.magic.gds
string GDS_START 23756
<< end >>

