magic
tech gf180mcuC
magscale 1 5
timestamp 1669966707
<< obsm1 >>
rect 672 855 109312 78833
<< metal2 >>
rect 336 79600 392 79900
rect 1344 79600 1400 79900
rect 2016 79600 2072 79900
rect 3024 79600 3080 79900
rect 4032 79600 4088 79900
rect 5040 79600 5096 79900
rect 5712 79600 5768 79900
rect 6720 79600 6776 79900
rect 7728 79600 7784 79900
rect 8400 79600 8456 79900
rect 9408 79600 9464 79900
rect 10416 79600 10472 79900
rect 11424 79600 11480 79900
rect 12096 79600 12152 79900
rect 13104 79600 13160 79900
rect 14112 79600 14168 79900
rect 14784 79600 14840 79900
rect 15792 79600 15848 79900
rect 16800 79600 16856 79900
rect 17808 79600 17864 79900
rect 18480 79600 18536 79900
rect 19488 79600 19544 79900
rect 20496 79600 20552 79900
rect 21504 79600 21560 79900
rect 22176 79600 22232 79900
rect 23184 79600 23240 79900
rect 24192 79600 24248 79900
rect 24864 79600 24920 79900
rect 25872 79600 25928 79900
rect 26880 79600 26936 79900
rect 27888 79600 27944 79900
rect 28560 79600 28616 79900
rect 29568 79600 29624 79900
rect 30576 79600 30632 79900
rect 31248 79600 31304 79900
rect 32256 79600 32312 79900
rect 33264 79600 33320 79900
rect 34272 79600 34328 79900
rect 34944 79600 35000 79900
rect 35952 79600 36008 79900
rect 36960 79600 37016 79900
rect 37968 79600 38024 79900
rect 38640 79600 38696 79900
rect 39648 79600 39704 79900
rect 40656 79600 40712 79900
rect 41328 79600 41384 79900
rect 42336 79600 42392 79900
rect 43344 79600 43400 79900
rect 44352 79600 44408 79900
rect 45024 79600 45080 79900
rect 46032 79600 46088 79900
rect 47040 79600 47096 79900
rect 47712 79600 47768 79900
rect 48720 79600 48776 79900
rect 49728 79600 49784 79900
rect 50736 79600 50792 79900
rect 51408 79600 51464 79900
rect 52416 79600 52472 79900
rect 53424 79600 53480 79900
rect 54432 79600 54488 79900
rect 55104 79600 55160 79900
rect 56112 79600 56168 79900
rect 57120 79600 57176 79900
rect 57792 79600 57848 79900
rect 58800 79600 58856 79900
rect 59808 79600 59864 79900
rect 60816 79600 60872 79900
rect 61488 79600 61544 79900
rect 62496 79600 62552 79900
rect 63504 79600 63560 79900
rect 64176 79600 64232 79900
rect 65184 79600 65240 79900
rect 66192 79600 66248 79900
rect 67200 79600 67256 79900
rect 67872 79600 67928 79900
rect 68880 79600 68936 79900
rect 69888 79600 69944 79900
rect 70560 79600 70616 79900
rect 71568 79600 71624 79900
rect 72576 79600 72632 79900
rect 73584 79600 73640 79900
rect 74256 79600 74312 79900
rect 75264 79600 75320 79900
rect 76272 79600 76328 79900
rect 77280 79600 77336 79900
rect 77952 79600 78008 79900
rect 78960 79600 79016 79900
rect 79968 79600 80024 79900
rect 80640 79600 80696 79900
rect 81648 79600 81704 79900
rect 82656 79600 82712 79900
rect 83664 79600 83720 79900
rect 84336 79600 84392 79900
rect 85344 79600 85400 79900
rect 86352 79600 86408 79900
rect 87024 79600 87080 79900
rect 88032 79600 88088 79900
rect 89040 79600 89096 79900
rect 90048 79600 90104 79900
rect 90720 79600 90776 79900
rect 91728 79600 91784 79900
rect 92736 79600 92792 79900
rect 93744 79600 93800 79900
rect 94416 79600 94472 79900
rect 95424 79600 95480 79900
rect 96432 79600 96488 79900
rect 97104 79600 97160 79900
rect 98112 79600 98168 79900
rect 99120 79600 99176 79900
rect 100128 79600 100184 79900
rect 100800 79600 100856 79900
rect 101808 79600 101864 79900
rect 102816 79600 102872 79900
rect 103488 79600 103544 79900
rect 104496 79600 104552 79900
rect 105504 79600 105560 79900
rect 106512 79600 106568 79900
rect 107184 79600 107240 79900
rect 108192 79600 108248 79900
rect 109200 79600 109256 79900
rect 109872 79600 109928 79900
rect 0 100 56 400
rect 672 100 728 400
rect 1680 100 1736 400
rect 2688 100 2744 400
rect 3360 100 3416 400
rect 4368 100 4424 400
rect 5376 100 5432 400
rect 6384 100 6440 400
rect 7056 100 7112 400
rect 8064 100 8120 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10752 100 10808 400
rect 11760 100 11816 400
rect 12768 100 12824 400
rect 13440 100 13496 400
rect 14448 100 14504 400
rect 15456 100 15512 400
rect 16128 100 16184 400
rect 17136 100 17192 400
rect 18144 100 18200 400
rect 19152 100 19208 400
rect 19824 100 19880 400
rect 20832 100 20888 400
rect 21840 100 21896 400
rect 22848 100 22904 400
rect 23520 100 23576 400
rect 24528 100 24584 400
rect 25536 100 25592 400
rect 26208 100 26264 400
rect 27216 100 27272 400
rect 28224 100 28280 400
rect 29232 100 29288 400
rect 29904 100 29960 400
rect 30912 100 30968 400
rect 31920 100 31976 400
rect 32592 100 32648 400
rect 33600 100 33656 400
rect 34608 100 34664 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 37296 100 37352 400
rect 38304 100 38360 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40992 100 41048 400
rect 42000 100 42056 400
rect 42672 100 42728 400
rect 43680 100 43736 400
rect 44688 100 44744 400
rect 45696 100 45752 400
rect 46368 100 46424 400
rect 47376 100 47432 400
rect 48384 100 48440 400
rect 49056 100 49112 400
rect 50064 100 50120 400
rect 51072 100 51128 400
rect 52080 100 52136 400
rect 52752 100 52808 400
rect 53760 100 53816 400
rect 54768 100 54824 400
rect 55440 100 55496 400
rect 56448 100 56504 400
rect 57456 100 57512 400
rect 58464 100 58520 400
rect 59136 100 59192 400
rect 60144 100 60200 400
rect 61152 100 61208 400
rect 62160 100 62216 400
rect 62832 100 62888 400
rect 63840 100 63896 400
rect 64848 100 64904 400
rect 65520 100 65576 400
rect 66528 100 66584 400
rect 67536 100 67592 400
rect 68544 100 68600 400
rect 69216 100 69272 400
rect 70224 100 70280 400
rect 71232 100 71288 400
rect 71904 100 71960 400
rect 72912 100 72968 400
rect 73920 100 73976 400
rect 74928 100 74984 400
rect 75600 100 75656 400
rect 76608 100 76664 400
rect 77616 100 77672 400
rect 78624 100 78680 400
rect 79296 100 79352 400
rect 80304 100 80360 400
rect 81312 100 81368 400
rect 81984 100 82040 400
rect 82992 100 83048 400
rect 84000 100 84056 400
rect 85008 100 85064 400
rect 85680 100 85736 400
rect 86688 100 86744 400
rect 87696 100 87752 400
rect 88368 100 88424 400
rect 89376 100 89432 400
rect 90384 100 90440 400
rect 91392 100 91448 400
rect 92064 100 92120 400
rect 93072 100 93128 400
rect 94080 100 94136 400
rect 95088 100 95144 400
rect 95760 100 95816 400
rect 96768 100 96824 400
rect 97776 100 97832 400
rect 98448 100 98504 400
rect 99456 100 99512 400
rect 100464 100 100520 400
rect 101472 100 101528 400
rect 102144 100 102200 400
rect 103152 100 103208 400
rect 104160 100 104216 400
rect 104832 100 104888 400
rect 105840 100 105896 400
rect 106848 100 106904 400
rect 107856 100 107912 400
rect 108528 100 108584 400
rect 109536 100 109592 400
<< obsm2 >>
rect 14 79570 306 79600
rect 422 79570 1314 79600
rect 1430 79570 1986 79600
rect 2102 79570 2994 79600
rect 3110 79570 4002 79600
rect 4118 79570 5010 79600
rect 5126 79570 5682 79600
rect 5798 79570 6690 79600
rect 6806 79570 7698 79600
rect 7814 79570 8370 79600
rect 8486 79570 9378 79600
rect 9494 79570 10386 79600
rect 10502 79570 11394 79600
rect 11510 79570 12066 79600
rect 12182 79570 13074 79600
rect 13190 79570 14082 79600
rect 14198 79570 14754 79600
rect 14870 79570 15762 79600
rect 15878 79570 16770 79600
rect 16886 79570 17778 79600
rect 17894 79570 18450 79600
rect 18566 79570 19458 79600
rect 19574 79570 20466 79600
rect 20582 79570 21474 79600
rect 21590 79570 22146 79600
rect 22262 79570 23154 79600
rect 23270 79570 24162 79600
rect 24278 79570 24834 79600
rect 24950 79570 25842 79600
rect 25958 79570 26850 79600
rect 26966 79570 27858 79600
rect 27974 79570 28530 79600
rect 28646 79570 29538 79600
rect 29654 79570 30546 79600
rect 30662 79570 31218 79600
rect 31334 79570 32226 79600
rect 32342 79570 33234 79600
rect 33350 79570 34242 79600
rect 34358 79570 34914 79600
rect 35030 79570 35922 79600
rect 36038 79570 36930 79600
rect 37046 79570 37938 79600
rect 38054 79570 38610 79600
rect 38726 79570 39618 79600
rect 39734 79570 40626 79600
rect 40742 79570 41298 79600
rect 41414 79570 42306 79600
rect 42422 79570 43314 79600
rect 43430 79570 44322 79600
rect 44438 79570 44994 79600
rect 45110 79570 46002 79600
rect 46118 79570 47010 79600
rect 47126 79570 47682 79600
rect 47798 79570 48690 79600
rect 48806 79570 49698 79600
rect 49814 79570 50706 79600
rect 50822 79570 51378 79600
rect 51494 79570 52386 79600
rect 52502 79570 53394 79600
rect 53510 79570 54402 79600
rect 54518 79570 55074 79600
rect 55190 79570 56082 79600
rect 56198 79570 57090 79600
rect 57206 79570 57762 79600
rect 57878 79570 58770 79600
rect 58886 79570 59778 79600
rect 59894 79570 60786 79600
rect 60902 79570 61458 79600
rect 61574 79570 62466 79600
rect 62582 79570 63474 79600
rect 63590 79570 64146 79600
rect 64262 79570 65154 79600
rect 65270 79570 66162 79600
rect 66278 79570 67170 79600
rect 67286 79570 67842 79600
rect 67958 79570 68850 79600
rect 68966 79570 69858 79600
rect 69974 79570 70530 79600
rect 70646 79570 71538 79600
rect 71654 79570 72546 79600
rect 72662 79570 73554 79600
rect 73670 79570 74226 79600
rect 74342 79570 75234 79600
rect 75350 79570 76242 79600
rect 76358 79570 77250 79600
rect 77366 79570 77922 79600
rect 78038 79570 78930 79600
rect 79046 79570 79938 79600
rect 80054 79570 80610 79600
rect 80726 79570 81618 79600
rect 81734 79570 82626 79600
rect 82742 79570 83634 79600
rect 83750 79570 84306 79600
rect 84422 79570 85314 79600
rect 85430 79570 86322 79600
rect 86438 79570 86994 79600
rect 87110 79570 88002 79600
rect 88118 79570 89010 79600
rect 89126 79570 90018 79600
rect 90134 79570 90690 79600
rect 90806 79570 91698 79600
rect 91814 79570 92706 79600
rect 92822 79570 93714 79600
rect 93830 79570 94386 79600
rect 94502 79570 95394 79600
rect 95510 79570 96402 79600
rect 96518 79570 97074 79600
rect 97190 79570 98082 79600
rect 98198 79570 99090 79600
rect 99206 79570 100098 79600
rect 100214 79570 100770 79600
rect 100886 79570 101778 79600
rect 101894 79570 102786 79600
rect 102902 79570 103458 79600
rect 103574 79570 104466 79600
rect 104582 79570 105474 79600
rect 105590 79570 106482 79600
rect 106598 79570 107154 79600
rect 107270 79570 108162 79600
rect 108278 79570 109074 79600
rect 14 430 109074 79570
rect 86 400 642 430
rect 758 400 1650 430
rect 1766 400 2658 430
rect 2774 400 3330 430
rect 3446 400 4338 430
rect 4454 400 5346 430
rect 5462 400 6354 430
rect 6470 400 7026 430
rect 7142 400 8034 430
rect 8150 400 9042 430
rect 9158 400 9714 430
rect 9830 400 10722 430
rect 10838 400 11730 430
rect 11846 400 12738 430
rect 12854 400 13410 430
rect 13526 400 14418 430
rect 14534 400 15426 430
rect 15542 400 16098 430
rect 16214 400 17106 430
rect 17222 400 18114 430
rect 18230 400 19122 430
rect 19238 400 19794 430
rect 19910 400 20802 430
rect 20918 400 21810 430
rect 21926 400 22818 430
rect 22934 400 23490 430
rect 23606 400 24498 430
rect 24614 400 25506 430
rect 25622 400 26178 430
rect 26294 400 27186 430
rect 27302 400 28194 430
rect 28310 400 29202 430
rect 29318 400 29874 430
rect 29990 400 30882 430
rect 30998 400 31890 430
rect 32006 400 32562 430
rect 32678 400 33570 430
rect 33686 400 34578 430
rect 34694 400 35586 430
rect 35702 400 36258 430
rect 36374 400 37266 430
rect 37382 400 38274 430
rect 38390 400 39282 430
rect 39398 400 39954 430
rect 40070 400 40962 430
rect 41078 400 41970 430
rect 42086 400 42642 430
rect 42758 400 43650 430
rect 43766 400 44658 430
rect 44774 400 45666 430
rect 45782 400 46338 430
rect 46454 400 47346 430
rect 47462 400 48354 430
rect 48470 400 49026 430
rect 49142 400 50034 430
rect 50150 400 51042 430
rect 51158 400 52050 430
rect 52166 400 52722 430
rect 52838 400 53730 430
rect 53846 400 54738 430
rect 54854 400 55410 430
rect 55526 400 56418 430
rect 56534 400 57426 430
rect 57542 400 58434 430
rect 58550 400 59106 430
rect 59222 400 60114 430
rect 60230 400 61122 430
rect 61238 400 62130 430
rect 62246 400 62802 430
rect 62918 400 63810 430
rect 63926 400 64818 430
rect 64934 400 65490 430
rect 65606 400 66498 430
rect 66614 400 67506 430
rect 67622 400 68514 430
rect 68630 400 69186 430
rect 69302 400 70194 430
rect 70310 400 71202 430
rect 71318 400 71874 430
rect 71990 400 72882 430
rect 72998 400 73890 430
rect 74006 400 74898 430
rect 75014 400 75570 430
rect 75686 400 76578 430
rect 76694 400 77586 430
rect 77702 400 78594 430
rect 78710 400 79266 430
rect 79382 400 80274 430
rect 80390 400 81282 430
rect 81398 400 81954 430
rect 82070 400 82962 430
rect 83078 400 83970 430
rect 84086 400 84978 430
rect 85094 400 85650 430
rect 85766 400 86658 430
rect 86774 400 87666 430
rect 87782 400 88338 430
rect 88454 400 89346 430
rect 89462 400 90354 430
rect 90470 400 91362 430
rect 91478 400 92034 430
rect 92150 400 93042 430
rect 93158 400 94050 430
rect 94166 400 95058 430
rect 95174 400 95730 430
rect 95846 400 96738 430
rect 96854 400 97746 430
rect 97862 400 98418 430
rect 98534 400 99426 430
rect 99542 400 100434 430
rect 100550 400 101442 430
rect 101558 400 102114 430
rect 102230 400 103122 430
rect 103238 400 104130 430
rect 104246 400 104802 430
rect 104918 400 105810 430
rect 105926 400 106818 430
rect 106934 400 107826 430
rect 107942 400 108498 430
rect 108614 400 109074 430
<< metal3 >>
rect 100 79296 400 79352
rect 109600 78960 109900 79016
rect 100 78624 400 78680
rect 109600 77952 109900 78008
rect 100 77616 400 77672
rect 109600 76944 109900 77000
rect 100 76608 400 76664
rect 109600 76272 109900 76328
rect 100 75600 400 75656
rect 109600 75264 109900 75320
rect 100 74928 400 74984
rect 109600 74256 109900 74312
rect 100 73920 400 73976
rect 109600 73248 109900 73304
rect 100 72912 400 72968
rect 109600 72576 109900 72632
rect 100 71904 400 71960
rect 109600 71568 109900 71624
rect 100 71232 400 71288
rect 109600 70560 109900 70616
rect 100 70224 400 70280
rect 109600 69888 109900 69944
rect 100 69216 400 69272
rect 109600 68880 109900 68936
rect 100 68544 400 68600
rect 109600 67872 109900 67928
rect 100 67536 400 67592
rect 109600 66864 109900 66920
rect 100 66528 400 66584
rect 109600 66192 109900 66248
rect 100 65520 400 65576
rect 109600 65184 109900 65240
rect 100 64848 400 64904
rect 109600 64176 109900 64232
rect 100 63840 400 63896
rect 109600 63504 109900 63560
rect 100 62832 400 62888
rect 109600 62496 109900 62552
rect 100 62160 400 62216
rect 109600 61488 109900 61544
rect 100 61152 400 61208
rect 109600 60480 109900 60536
rect 100 60144 400 60200
rect 109600 59808 109900 59864
rect 100 59136 400 59192
rect 109600 58800 109900 58856
rect 100 58464 400 58520
rect 109600 57792 109900 57848
rect 100 57456 400 57512
rect 109600 56784 109900 56840
rect 100 56448 400 56504
rect 109600 56112 109900 56168
rect 100 55440 400 55496
rect 109600 55104 109900 55160
rect 100 54768 400 54824
rect 109600 54096 109900 54152
rect 100 53760 400 53816
rect 109600 53424 109900 53480
rect 100 52752 400 52808
rect 109600 52416 109900 52472
rect 100 52080 400 52136
rect 109600 51408 109900 51464
rect 100 51072 400 51128
rect 109600 50400 109900 50456
rect 100 50064 400 50120
rect 109600 49728 109900 49784
rect 100 49056 400 49112
rect 109600 48720 109900 48776
rect 100 48384 400 48440
rect 109600 47712 109900 47768
rect 100 47376 400 47432
rect 109600 47040 109900 47096
rect 100 46368 400 46424
rect 109600 46032 109900 46088
rect 100 45696 400 45752
rect 109600 45024 109900 45080
rect 100 44688 400 44744
rect 109600 44016 109900 44072
rect 100 43680 400 43736
rect 109600 43344 109900 43400
rect 100 42672 400 42728
rect 109600 42336 109900 42392
rect 100 42000 400 42056
rect 109600 41328 109900 41384
rect 100 40992 400 41048
rect 109600 40320 109900 40376
rect 100 39984 400 40040
rect 109600 39648 109900 39704
rect 100 39312 400 39368
rect 109600 38640 109900 38696
rect 100 38304 400 38360
rect 109600 37632 109900 37688
rect 100 37296 400 37352
rect 109600 36960 109900 37016
rect 100 36288 400 36344
rect 109600 35952 109900 36008
rect 100 35616 400 35672
rect 109600 34944 109900 35000
rect 100 34608 400 34664
rect 109600 33936 109900 33992
rect 100 33600 400 33656
rect 109600 33264 109900 33320
rect 100 32592 400 32648
rect 109600 32256 109900 32312
rect 100 31920 400 31976
rect 109600 31248 109900 31304
rect 100 30912 400 30968
rect 109600 30576 109900 30632
rect 100 29904 400 29960
rect 109600 29568 109900 29624
rect 100 29232 400 29288
rect 109600 28560 109900 28616
rect 100 28224 400 28280
rect 109600 27552 109900 27608
rect 100 27216 400 27272
rect 109600 26880 109900 26936
rect 100 26208 400 26264
rect 109600 25872 109900 25928
rect 100 25536 400 25592
rect 109600 24864 109900 24920
rect 100 24528 400 24584
rect 109600 24192 109900 24248
rect 100 23520 400 23576
rect 109600 23184 109900 23240
rect 100 22848 400 22904
rect 109600 22176 109900 22232
rect 100 21840 400 21896
rect 109600 21168 109900 21224
rect 100 20832 400 20888
rect 109600 20496 109900 20552
rect 100 19824 400 19880
rect 109600 19488 109900 19544
rect 100 19152 400 19208
rect 109600 18480 109900 18536
rect 100 18144 400 18200
rect 109600 17472 109900 17528
rect 100 17136 400 17192
rect 109600 16800 109900 16856
rect 100 16128 400 16184
rect 109600 15792 109900 15848
rect 100 15456 400 15512
rect 109600 14784 109900 14840
rect 100 14448 400 14504
rect 109600 14112 109900 14168
rect 100 13440 400 13496
rect 109600 13104 109900 13160
rect 100 12768 400 12824
rect 109600 12096 109900 12152
rect 100 11760 400 11816
rect 109600 11088 109900 11144
rect 100 10752 400 10808
rect 109600 10416 109900 10472
rect 100 9744 400 9800
rect 109600 9408 109900 9464
rect 100 9072 400 9128
rect 109600 8400 109900 8456
rect 100 8064 400 8120
rect 109600 7728 109900 7784
rect 100 7056 400 7112
rect 109600 6720 109900 6776
rect 100 6384 400 6440
rect 109600 5712 109900 5768
rect 100 5376 400 5432
rect 109600 4704 109900 4760
rect 100 4368 400 4424
rect 109600 4032 109900 4088
rect 100 3360 400 3416
rect 109600 3024 109900 3080
rect 100 2688 400 2744
rect 109600 2016 109900 2072
rect 100 1680 400 1736
rect 109600 1008 109900 1064
rect 100 672 400 728
rect 109600 336 109900 392
<< obsm3 >>
rect 9 78038 109970 78414
rect 9 77922 109570 78038
rect 109930 77922 109970 78038
rect 9 77702 109970 77922
rect 9 77586 70 77702
rect 430 77586 109970 77702
rect 9 77030 109970 77586
rect 9 76914 109570 77030
rect 109930 76914 109970 77030
rect 9 76694 109970 76914
rect 9 76578 70 76694
rect 430 76578 109970 76694
rect 9 76358 109970 76578
rect 9 76242 109570 76358
rect 109930 76242 109970 76358
rect 9 75686 109970 76242
rect 9 75570 70 75686
rect 430 75570 109970 75686
rect 9 75350 109970 75570
rect 9 75234 109570 75350
rect 109930 75234 109970 75350
rect 9 75014 109970 75234
rect 9 74898 70 75014
rect 430 74898 109970 75014
rect 9 74342 109970 74898
rect 9 74226 109570 74342
rect 109930 74226 109970 74342
rect 9 74006 109970 74226
rect 9 73890 70 74006
rect 430 73890 109970 74006
rect 9 73334 109970 73890
rect 9 73218 109570 73334
rect 109930 73218 109970 73334
rect 9 72998 109970 73218
rect 9 72882 70 72998
rect 430 72882 109970 72998
rect 9 72662 109970 72882
rect 9 72546 109570 72662
rect 109930 72546 109970 72662
rect 9 71990 109970 72546
rect 9 71874 70 71990
rect 430 71874 109970 71990
rect 9 71654 109970 71874
rect 9 71538 109570 71654
rect 109930 71538 109970 71654
rect 9 71318 109970 71538
rect 9 71202 70 71318
rect 430 71202 109970 71318
rect 9 70646 109970 71202
rect 9 70530 109570 70646
rect 109930 70530 109970 70646
rect 9 70310 109970 70530
rect 9 70194 70 70310
rect 430 70194 109970 70310
rect 9 69974 109970 70194
rect 9 69858 109570 69974
rect 109930 69858 109970 69974
rect 9 69302 109970 69858
rect 9 69186 70 69302
rect 430 69186 109970 69302
rect 9 68966 109970 69186
rect 9 68850 109570 68966
rect 109930 68850 109970 68966
rect 9 68630 109970 68850
rect 9 68514 70 68630
rect 430 68514 109970 68630
rect 9 67958 109970 68514
rect 9 67842 109570 67958
rect 109930 67842 109970 67958
rect 9 67622 109970 67842
rect 9 67506 70 67622
rect 430 67506 109970 67622
rect 9 66950 109970 67506
rect 9 66834 109570 66950
rect 109930 66834 109970 66950
rect 9 66614 109970 66834
rect 9 66498 70 66614
rect 430 66498 109970 66614
rect 9 66278 109970 66498
rect 9 66162 109570 66278
rect 109930 66162 109970 66278
rect 9 65606 109970 66162
rect 9 65490 70 65606
rect 430 65490 109970 65606
rect 9 65270 109970 65490
rect 9 65154 109570 65270
rect 109930 65154 109970 65270
rect 9 64934 109970 65154
rect 9 64818 70 64934
rect 430 64818 109970 64934
rect 9 64262 109970 64818
rect 9 64146 109570 64262
rect 109930 64146 109970 64262
rect 9 63926 109970 64146
rect 9 63810 70 63926
rect 430 63810 109970 63926
rect 9 63590 109970 63810
rect 9 63474 109570 63590
rect 109930 63474 109970 63590
rect 9 62918 109970 63474
rect 9 62802 70 62918
rect 430 62802 109970 62918
rect 9 62582 109970 62802
rect 9 62466 109570 62582
rect 109930 62466 109970 62582
rect 9 62246 109970 62466
rect 9 62130 70 62246
rect 430 62130 109970 62246
rect 9 61574 109970 62130
rect 9 61458 109570 61574
rect 109930 61458 109970 61574
rect 9 61238 109970 61458
rect 9 61122 70 61238
rect 430 61122 109970 61238
rect 9 60566 109970 61122
rect 9 60450 109570 60566
rect 109930 60450 109970 60566
rect 9 60230 109970 60450
rect 9 60114 70 60230
rect 430 60114 109970 60230
rect 9 59894 109970 60114
rect 9 59778 109570 59894
rect 109930 59778 109970 59894
rect 9 59222 109970 59778
rect 9 59106 70 59222
rect 430 59106 109970 59222
rect 9 58886 109970 59106
rect 9 58770 109570 58886
rect 109930 58770 109970 58886
rect 9 58550 109970 58770
rect 9 58434 70 58550
rect 430 58434 109970 58550
rect 9 57878 109970 58434
rect 9 57762 109570 57878
rect 109930 57762 109970 57878
rect 9 57542 109970 57762
rect 9 57426 70 57542
rect 430 57426 109970 57542
rect 9 56870 109970 57426
rect 9 56754 109570 56870
rect 109930 56754 109970 56870
rect 9 56534 109970 56754
rect 9 56418 70 56534
rect 430 56418 109970 56534
rect 9 56198 109970 56418
rect 9 56082 109570 56198
rect 109930 56082 109970 56198
rect 9 55526 109970 56082
rect 9 55410 70 55526
rect 430 55410 109970 55526
rect 9 55190 109970 55410
rect 9 55074 109570 55190
rect 109930 55074 109970 55190
rect 9 54854 109970 55074
rect 9 54738 70 54854
rect 430 54738 109970 54854
rect 9 54182 109970 54738
rect 9 54066 109570 54182
rect 109930 54066 109970 54182
rect 9 53846 109970 54066
rect 9 53730 70 53846
rect 430 53730 109970 53846
rect 9 53510 109970 53730
rect 9 53394 109570 53510
rect 109930 53394 109970 53510
rect 9 52838 109970 53394
rect 9 52722 70 52838
rect 430 52722 109970 52838
rect 9 52502 109970 52722
rect 9 52386 109570 52502
rect 109930 52386 109970 52502
rect 9 52166 109970 52386
rect 9 52050 70 52166
rect 430 52050 109970 52166
rect 9 51494 109970 52050
rect 9 51378 109570 51494
rect 109930 51378 109970 51494
rect 9 51158 109970 51378
rect 9 51042 70 51158
rect 430 51042 109970 51158
rect 9 50486 109970 51042
rect 9 50370 109570 50486
rect 109930 50370 109970 50486
rect 9 50150 109970 50370
rect 9 50034 70 50150
rect 430 50034 109970 50150
rect 9 49814 109970 50034
rect 9 49698 109570 49814
rect 109930 49698 109970 49814
rect 9 49142 109970 49698
rect 9 49026 70 49142
rect 430 49026 109970 49142
rect 9 48806 109970 49026
rect 9 48690 109570 48806
rect 109930 48690 109970 48806
rect 9 48470 109970 48690
rect 9 48354 70 48470
rect 430 48354 109970 48470
rect 9 47798 109970 48354
rect 9 47682 109570 47798
rect 109930 47682 109970 47798
rect 9 47462 109970 47682
rect 9 47346 70 47462
rect 430 47346 109970 47462
rect 9 47126 109970 47346
rect 9 47010 109570 47126
rect 109930 47010 109970 47126
rect 9 46454 109970 47010
rect 9 46338 70 46454
rect 430 46338 109970 46454
rect 9 46118 109970 46338
rect 9 46002 109570 46118
rect 109930 46002 109970 46118
rect 9 45782 109970 46002
rect 9 45666 70 45782
rect 430 45666 109970 45782
rect 9 45110 109970 45666
rect 9 44994 109570 45110
rect 109930 44994 109970 45110
rect 9 44774 109970 44994
rect 9 44658 70 44774
rect 430 44658 109970 44774
rect 9 44102 109970 44658
rect 9 43986 109570 44102
rect 109930 43986 109970 44102
rect 9 43766 109970 43986
rect 9 43650 70 43766
rect 430 43650 109970 43766
rect 9 43430 109970 43650
rect 9 43314 109570 43430
rect 109930 43314 109970 43430
rect 9 42758 109970 43314
rect 9 42642 70 42758
rect 430 42642 109970 42758
rect 9 42422 109970 42642
rect 9 42306 109570 42422
rect 109930 42306 109970 42422
rect 9 42086 109970 42306
rect 9 41970 70 42086
rect 430 41970 109970 42086
rect 9 41414 109970 41970
rect 9 41298 109570 41414
rect 109930 41298 109970 41414
rect 9 41078 109970 41298
rect 9 40962 70 41078
rect 430 40962 109970 41078
rect 9 40406 109970 40962
rect 9 40290 109570 40406
rect 109930 40290 109970 40406
rect 9 40070 109970 40290
rect 9 39954 70 40070
rect 430 39954 109970 40070
rect 9 39734 109970 39954
rect 9 39618 109570 39734
rect 109930 39618 109970 39734
rect 9 39398 109970 39618
rect 9 39282 70 39398
rect 430 39282 109970 39398
rect 9 38726 109970 39282
rect 9 38610 109570 38726
rect 109930 38610 109970 38726
rect 9 38390 109970 38610
rect 9 38274 70 38390
rect 430 38274 109970 38390
rect 9 37718 109970 38274
rect 9 37602 109570 37718
rect 109930 37602 109970 37718
rect 9 37382 109970 37602
rect 9 37266 70 37382
rect 430 37266 109970 37382
rect 9 37046 109970 37266
rect 9 36930 109570 37046
rect 109930 36930 109970 37046
rect 9 36374 109970 36930
rect 9 36258 70 36374
rect 430 36258 109970 36374
rect 9 36038 109970 36258
rect 9 35922 109570 36038
rect 109930 35922 109970 36038
rect 9 35702 109970 35922
rect 9 35586 70 35702
rect 430 35586 109970 35702
rect 9 35030 109970 35586
rect 9 34914 109570 35030
rect 109930 34914 109970 35030
rect 9 34694 109970 34914
rect 9 34578 70 34694
rect 430 34578 109970 34694
rect 9 34022 109970 34578
rect 9 33906 109570 34022
rect 109930 33906 109970 34022
rect 9 33686 109970 33906
rect 9 33570 70 33686
rect 430 33570 109970 33686
rect 9 33350 109970 33570
rect 9 33234 109570 33350
rect 109930 33234 109970 33350
rect 9 32678 109970 33234
rect 9 32562 70 32678
rect 430 32562 109970 32678
rect 9 32342 109970 32562
rect 9 32226 109570 32342
rect 109930 32226 109970 32342
rect 9 32006 109970 32226
rect 9 31890 70 32006
rect 430 31890 109970 32006
rect 9 31334 109970 31890
rect 9 31218 109570 31334
rect 109930 31218 109970 31334
rect 9 30998 109970 31218
rect 9 30882 70 30998
rect 430 30882 109970 30998
rect 9 30662 109970 30882
rect 9 30546 109570 30662
rect 109930 30546 109970 30662
rect 9 29990 109970 30546
rect 9 29874 70 29990
rect 430 29874 109970 29990
rect 9 29654 109970 29874
rect 9 29538 109570 29654
rect 109930 29538 109970 29654
rect 9 29318 109970 29538
rect 9 29202 70 29318
rect 430 29202 109970 29318
rect 9 28646 109970 29202
rect 9 28530 109570 28646
rect 109930 28530 109970 28646
rect 9 28310 109970 28530
rect 9 28194 70 28310
rect 430 28194 109970 28310
rect 9 27638 109970 28194
rect 9 27522 109570 27638
rect 109930 27522 109970 27638
rect 9 27302 109970 27522
rect 9 27186 70 27302
rect 430 27186 109970 27302
rect 9 26966 109970 27186
rect 9 26850 109570 26966
rect 109930 26850 109970 26966
rect 9 26294 109970 26850
rect 9 26178 70 26294
rect 430 26178 109970 26294
rect 9 25958 109970 26178
rect 9 25842 109570 25958
rect 109930 25842 109970 25958
rect 9 25622 109970 25842
rect 9 25506 70 25622
rect 430 25506 109970 25622
rect 9 24950 109970 25506
rect 9 24834 109570 24950
rect 109930 24834 109970 24950
rect 9 24614 109970 24834
rect 9 24498 70 24614
rect 430 24498 109970 24614
rect 9 24278 109970 24498
rect 9 24162 109570 24278
rect 109930 24162 109970 24278
rect 9 23606 109970 24162
rect 9 23490 70 23606
rect 430 23490 109970 23606
rect 9 23270 109970 23490
rect 9 23154 109570 23270
rect 109930 23154 109970 23270
rect 9 22934 109970 23154
rect 9 22818 70 22934
rect 430 22818 109970 22934
rect 9 22262 109970 22818
rect 9 22146 109570 22262
rect 109930 22146 109970 22262
rect 9 21926 109970 22146
rect 9 21810 70 21926
rect 430 21810 109970 21926
rect 9 21254 109970 21810
rect 9 21138 109570 21254
rect 109930 21138 109970 21254
rect 9 20918 109970 21138
rect 9 20802 70 20918
rect 430 20802 109970 20918
rect 9 20582 109970 20802
rect 9 20466 109570 20582
rect 109930 20466 109970 20582
rect 9 19910 109970 20466
rect 9 19794 70 19910
rect 430 19794 109970 19910
rect 9 19574 109970 19794
rect 9 19458 109570 19574
rect 109930 19458 109970 19574
rect 9 19238 109970 19458
rect 9 19122 70 19238
rect 430 19122 109970 19238
rect 9 18566 109970 19122
rect 9 18450 109570 18566
rect 109930 18450 109970 18566
rect 9 18230 109970 18450
rect 9 18114 70 18230
rect 430 18114 109970 18230
rect 9 17558 109970 18114
rect 9 17442 109570 17558
rect 109930 17442 109970 17558
rect 9 17222 109970 17442
rect 9 17106 70 17222
rect 430 17106 109970 17222
rect 9 16886 109970 17106
rect 9 16770 109570 16886
rect 109930 16770 109970 16886
rect 9 16214 109970 16770
rect 9 16098 70 16214
rect 430 16098 109970 16214
rect 9 15878 109970 16098
rect 9 15762 109570 15878
rect 109930 15762 109970 15878
rect 9 15542 109970 15762
rect 9 15426 70 15542
rect 430 15426 109970 15542
rect 9 14870 109970 15426
rect 9 14754 109570 14870
rect 109930 14754 109970 14870
rect 9 14534 109970 14754
rect 9 14418 70 14534
rect 430 14418 109970 14534
rect 9 14198 109970 14418
rect 9 14082 109570 14198
rect 109930 14082 109970 14198
rect 9 13526 109970 14082
rect 9 13410 70 13526
rect 430 13410 109970 13526
rect 9 13190 109970 13410
rect 9 13074 109570 13190
rect 109930 13074 109970 13190
rect 9 12854 109970 13074
rect 9 12738 70 12854
rect 430 12738 109970 12854
rect 9 12182 109970 12738
rect 9 12066 109570 12182
rect 109930 12066 109970 12182
rect 9 11846 109970 12066
rect 9 11730 70 11846
rect 430 11730 109970 11846
rect 9 11174 109970 11730
rect 9 11058 109570 11174
rect 109930 11058 109970 11174
rect 9 10838 109970 11058
rect 9 10722 70 10838
rect 430 10722 109970 10838
rect 9 10502 109970 10722
rect 9 10386 109570 10502
rect 109930 10386 109970 10502
rect 9 9830 109970 10386
rect 9 9714 70 9830
rect 430 9714 109970 9830
rect 9 9494 109970 9714
rect 9 9378 109570 9494
rect 109930 9378 109970 9494
rect 9 9158 109970 9378
rect 9 9042 70 9158
rect 430 9042 109970 9158
rect 9 8486 109970 9042
rect 9 8370 109570 8486
rect 109930 8370 109970 8486
rect 9 8150 109970 8370
rect 9 8034 70 8150
rect 430 8034 109970 8150
rect 9 7814 109970 8034
rect 9 7698 109570 7814
rect 109930 7698 109970 7814
rect 9 7142 109970 7698
rect 9 7026 70 7142
rect 430 7026 109970 7142
rect 9 6806 109970 7026
rect 9 6690 109570 6806
rect 109930 6690 109970 6806
rect 9 6470 109970 6690
rect 9 6354 70 6470
rect 430 6354 109970 6470
rect 9 5798 109970 6354
rect 9 5682 109570 5798
rect 109930 5682 109970 5798
rect 9 5462 109970 5682
rect 9 5346 70 5462
rect 430 5346 109970 5462
rect 9 4790 109970 5346
rect 9 4674 109570 4790
rect 109930 4674 109970 4790
rect 9 4454 109970 4674
rect 9 4338 70 4454
rect 430 4338 109970 4454
rect 9 4118 109970 4338
rect 9 4002 109570 4118
rect 109930 4002 109970 4118
rect 9 3446 109970 4002
rect 9 3330 70 3446
rect 430 3330 109970 3446
rect 9 3110 109970 3330
rect 9 2994 109570 3110
rect 109930 2994 109970 3110
rect 9 2774 109970 2994
rect 9 2658 70 2774
rect 430 2658 109970 2774
rect 9 2102 109970 2658
rect 9 1986 109570 2102
rect 109930 1986 109970 2102
rect 9 1766 109970 1986
rect 9 1650 70 1766
rect 430 1650 109970 1766
rect 9 1094 109970 1650
rect 9 978 109570 1094
rect 109930 978 109970 1094
rect 9 758 109970 978
rect 9 642 70 758
rect 430 642 109970 758
rect 9 422 109970 642
rect 9 350 109570 422
rect 109930 350 109970 422
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
rect 86704 1538 86864 78430
rect 94384 1538 94544 78430
rect 102064 1538 102224 78430
<< labels >>
rlabel metal3 s 100 65520 400 65576 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 32592 400 32648 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 57456 400 57512 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 65184 79600 65240 79900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 109600 4032 109900 4088 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 109600 74256 109900 74312 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 78960 79600 79016 79900 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 93072 100 93128 400 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 26880 79600 26936 79900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 90720 79600 90776 79900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 109872 79600 109928 79900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 109600 66864 109900 66920 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 78624 100 78680 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 12768 100 12824 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 79296 400 79352 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 64848 400 64904 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 73920 400 73976 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 59136 400 59192 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 109600 78960 109900 79016 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 62160 100 62216 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 39984 400 40040 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 80304 100 80360 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 9744 400 9800 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 5040 79600 5096 79900 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 100128 79600 100184 79900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 109600 68880 109900 68936 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 109600 56784 109900 56840 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 109600 77952 109900 78008 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 109600 27552 109900 27608 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 18144 400 18200 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 109600 3024 109900 3080 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 92736 79600 92792 79900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 109600 51408 109900 51464 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 109600 46032 109900 46088 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 18480 79600 18536 79900 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 58464 100 58520 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 24528 400 24584 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 86688 100 86744 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 75264 79600 75320 79900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 27216 100 27272 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 9072 100 9128 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 19488 79600 19544 79900 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 48720 79600 48776 79900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 40656 79600 40712 79900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 69888 79600 69944 79900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 81312 100 81368 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 109600 9408 109900 9464 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 107184 79600 107240 79900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 27216 400 27272 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 13440 400 13496 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 6720 79600 6776 79900 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 79296 100 79352 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 16800 79600 16856 79900 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 109600 33264 109900 33320 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 109600 21168 109900 21224 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 89376 100 89432 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 29232 400 29288 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 98112 79600 98168 79900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 109600 336 109900 392 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 77616 400 77672 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 109600 70560 109900 70616 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 67872 79600 67928 79900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 109600 23184 109900 23240 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 71232 400 71288 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 12768 400 12824 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 84336 79600 84392 79900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 74928 400 74984 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 60816 79600 60872 79900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 109600 76944 109900 77000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 30576 79600 30632 79900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 44352 79600 44408 79900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 61152 100 61208 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 108192 79600 108248 79900 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 14784 79600 14840 79900 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 70224 400 70280 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 109600 64176 109900 64232 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 10752 100 10808 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 88368 100 88424 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 35952 79600 36008 79900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6384 100 6440 400 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 104160 100 104216 400 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 62832 400 62888 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 109600 5712 109900 5768 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 35616 400 35672 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 82992 100 83048 400 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 97776 100 97832 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 39984 100 40040 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 31920 100 31976 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 81648 79600 81704 79900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 64848 100 64904 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 109600 18480 109900 18536 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 101808 79600 101864 79900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 33600 100 33656 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 74256 79600 74312 79900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 34608 400 34664 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 62832 100 62888 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56448 100 56504 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 22848 100 22904 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 4368 400 4424 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 58800 79600 58856 79900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 43680 100 43736 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 55104 79600 55160 79900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 17136 400 17192 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 53760 400 53816 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 69216 100 69272 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 24528 100 24584 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 48384 400 48440 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 109600 73248 109900 73304 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 109600 26880 109900 26936 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 29232 100 29288 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 53424 79600 53480 79900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 3024 79600 3080 79900 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 109600 53424 109900 53480 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 24192 79600 24248 79900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 109536 100 109592 400 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 62496 79600 62552 79900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 36960 79600 37016 79900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 109600 4704 109900 4760 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 71904 400 71960 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 42000 400 42056 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 109600 56112 109900 56168 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 63504 79600 63560 79900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 34944 79600 35000 79900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 73584 79600 73640 79900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 5712 79600 5768 79900 6 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 9408 79600 9464 79900 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 109600 8400 109900 8456 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 57120 79600 57176 79900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 7056 400 7112 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 95424 79600 95480 79900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 38304 400 38360 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 63840 400 63896 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 22176 79600 22232 79900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 4032 79600 4088 79900 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 67536 100 67592 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 13104 79600 13160 79900 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 42672 100 42728 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 67200 79600 67256 79900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 109600 36960 109900 37016 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 32592 100 32648 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 45696 100 45752 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 31920 400 31976 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 104496 79600 104552 79900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 95760 100 95816 400 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 30912 100 30968 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 109600 54096 109900 54152 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 59136 100 59192 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 59808 79600 59864 79900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 51408 79600 51464 79900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 23184 79600 23240 79900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 52416 79600 52472 79900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 44688 100 44744 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 109600 16800 109900 16856 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 89040 79600 89096 79900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 82656 79600 82712 79900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 25536 400 25592 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 17808 79600 17864 79900 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 34608 100 34664 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 109600 71568 109900 71624 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 16128 100 16184 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 109600 47712 109900 47768 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 2688 400 2744 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 55440 100 55496 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 39648 79600 39704 79900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 19152 100 19208 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 109600 19488 109900 19544 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 100800 79600 100856 79900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 97104 79600 97160 79900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 109600 35952 109900 36008 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 68544 400 68600 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 35616 100 35672 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 109600 24192 109900 24248 6 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 1344 79600 1400 79900 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 109600 37632 109900 37688 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 61488 79600 61544 79900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 109600 63504 109900 63560 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 50064 100 50120 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 109600 29568 109900 29624 6 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 108528 100 108584 400 6 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 14112 79600 14168 79900 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 109600 44016 109900 44072 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 28224 100 28280 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 42672 400 42728 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 51072 100 51128 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 12096 79600 12152 79900 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 72576 79600 72632 79900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 109600 60480 109900 60536 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 40992 100 41048 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 21840 400 21896 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 109600 28560 109900 28616 6 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 99456 100 99512 400 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 70560 79600 70616 79900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 109600 2016 109900 2072 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 46368 100 46424 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 66192 79600 66248 79900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 109600 61488 109900 61544 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 109600 22176 109900 22232 6 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 96768 100 96824 400 6 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 107856 100 107912 400 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 15456 400 15512 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 92064 100 92120 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 109600 14112 109900 14168 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 109600 65184 109900 65240 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 5376 100 5432 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 29568 79600 29624 79900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 28560 79600 28616 79900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 67536 400 67592 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 21840 100 21896 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 85680 100 85736 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 68880 79600 68936 79900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 47712 79600 47768 79900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 11424 79600 11480 79900 6 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 101472 100 101528 400 6 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 10416 79600 10472 79900 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 109600 49728 109900 49784 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 50736 79600 50792 79900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 109600 7728 109900 7784 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 87024 79600 87080 79900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 109600 50400 109900 50456 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 36288 400 36344 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 109600 41328 109900 41384 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 91728 79600 91784 79900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 25536 100 25592 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 81984 100 82040 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 102144 100 102200 400 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 109600 12096 109900 12152 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 106512 79600 106568 79900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 5376 400 5432 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 109600 30576 109900 30632 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 109600 20496 109900 20552 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 109600 52416 109900 52472 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 109600 38640 109900 38696 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 15792 79600 15848 79900 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 75600 400 75656 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 70224 100 70280 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 84000 100 84056 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 13440 100 13496 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 11760 400 11816 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 21504 79600 21560 79900 6 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 103152 100 103208 400 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 33264 79600 33320 79900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 55440 400 55496 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 54432 79600 54488 79900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 85344 79600 85400 79900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 26208 100 26264 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 109600 43344 109900 43400 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 85008 100 85064 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 34272 79600 34328 79900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 17136 100 17192 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 109600 75264 109900 75320 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 109200 79600 109256 79900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 109600 66192 109900 66248 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 56112 79600 56168 79900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 109600 62496 109900 62552 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 48384 100 48440 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 31248 79600 31304 79900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 27888 79600 27944 79900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 40992 400 41048 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 52080 400 52136 6 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 106848 100 106904 400 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 49728 79600 49784 79900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 60144 400 60200 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 93744 79600 93800 79900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 75600 100 75656 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 10752 400 10808 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 69216 400 69272 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 8400 79600 8456 79900 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 72912 100 72968 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 46032 79600 46088 79900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 94080 100 94136 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 109600 45024 109900 45080 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 51072 400 51128 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 109600 33936 109900 33992 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 71904 100 71960 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 99120 79600 99176 79900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 104832 100 104888 400 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 71568 79600 71624 79900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 87696 100 87752 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 46368 400 46424 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 11760 100 11816 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 109600 32256 109900 32312 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 22848 400 22904 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 109600 47040 109900 47096 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 23520 100 23576 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 90384 100 90440 400 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 42336 79600 42392 79900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 96432 79600 96488 79900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 109600 57792 109900 57848 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 38640 79600 38696 79900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 61152 400 61208 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 78430 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 78430 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 109600 1008 109900 1064 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 32256 79600 32312 79900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 109600 17472 109900 17528 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 77952 79600 78008 79900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 57792 79600 57848 79900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 54768 400 54824 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 8064 100 8120 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 52752 100 52808 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 9072 400 9128 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 109600 48720 109900 48776 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 60144 100 60200 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 109600 14784 109900 14840 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 91392 100 91448 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 6384 400 6440 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 103488 79600 103544 79900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 53760 100 53816 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 76608 100 76664 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 109600 6720 109900 6776 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 25872 79600 25928 79900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 16128 400 16184 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 47040 79600 47096 79900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 109600 40320 109900 40376 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 109600 76272 109900 76328 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 37296 100 37352 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 37296 400 37352 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 109600 24864 109900 24920 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 73920 100 73976 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 88032 79600 88088 79900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 71232 100 71288 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 23520 400 23576 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 4368 100 4424 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 95088 100 95144 400 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 109600 10416 109900 10472 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 45024 79600 45080 79900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 109600 67872 109900 67928 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 72912 400 72968 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 336 79600 392 79900 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 76608 400 76664 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 19824 400 19880 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 109600 34944 109900 35000 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 54768 100 54824 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 79968 79600 80024 79900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 102816 79600 102872 79900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 20496 79600 20552 79900 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 14448 100 14504 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 44688 400 44744 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 105504 79600 105560 79900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 109600 59808 109900 59864 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 109600 15792 109900 15848 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 65520 100 65576 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 94416 79600 94472 79900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 37968 79600 38024 79900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 29904 100 29960 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 109600 42336 109900 42392 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 77616 100 77672 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 109600 13104 109900 13160 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 98448 100 98504 400 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 15456 100 15512 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 47376 100 47432 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 109600 25872 109900 25928 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 90048 79600 90104 79900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 109600 69888 109900 69944 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 100464 100 100520 400 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 19152 400 19208 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 109600 39648 109900 39704 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1680 100 1736 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 109600 72576 109900 72632 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 86352 79600 86408 79900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 105840 100 105896 400 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 83664 79600 83720 79900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 26208 400 26264 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 29904 400 29960 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 63840 100 63896 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 74928 100 74984 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 45696 400 45752 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 2016 79600 2072 79900 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 41328 79600 41384 79900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 30912 400 30968 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 19824 100 19880 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 7056 100 7112 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 64176 79600 64232 79900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 43344 79600 43400 79900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 52080 100 52136 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 80640 79600 80696 79900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 109600 11088 109900 11144 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 62160 400 62216 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 109600 58800 109900 58856 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 20832 100 20888 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 36288 100 36344 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 8064 400 8120 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 109600 55104 109900 55160 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 57456 100 57512 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 77280 79600 77336 79900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 76272 79600 76328 79900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 7728 79600 7784 79900 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 24864 79600 24920 79900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 68544 100 68600 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 20832 400 20888 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 78624 400 78680 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 109600 31248 109900 31304 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3168290
string GDS_FILE /home/runner/work/tiny_user_project/tiny_user_project/openlane/tiny_user_project/runs/22_12_02_07_36/results/signoff/tiny_user_project.magic.gds
string GDS_START 48106
<< end >>

