magic
tech sky130A
magscale 1 2
timestamp 1662455659
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 179754 117552
<< metal2 >>
rect 32862 119200 32918 120000
rect 69570 119200 69626 120000
rect 106278 119200 106334 120000
rect 142986 119200 143042 120000
rect 179694 119200 179750 120000
rect 18 0 74 800
rect 36726 0 36782 800
rect 73434 0 73490 800
rect 110142 0 110198 800
rect 146850 0 146906 800
<< obsm2 >>
rect 1398 119144 32806 119354
rect 32974 119144 69514 119354
rect 69682 119144 106222 119354
rect 106390 119144 142930 119354
rect 143098 119144 179638 119354
rect 1398 856 179748 119144
rect 1398 800 36670 856
rect 36838 800 73378 856
rect 73546 800 110086 856
rect 110254 800 146794 856
rect 146962 800 179748 856
<< metal3 >>
rect 0 116288 800 116408
rect 179200 80928 180000 81048
rect 0 77528 800 77648
rect 179200 42168 180000 42288
rect 0 38768 800 38888
rect 179200 3408 180000 3528
<< obsm3 >>
rect 800 116488 179200 117537
rect 880 116208 179200 116488
rect 800 81128 179200 116208
rect 800 80848 179120 81128
rect 800 77728 179200 80848
rect 880 77448 179200 77728
rect 800 42368 179200 77448
rect 800 42088 179120 42368
rect 800 38968 179200 42088
rect 880 38688 179200 38968
rect 800 3608 179200 38688
rect 800 3328 179120 3608
rect 800 2143 179200 3328
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal3 s 179200 42168 180000 42288 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 32862 119200 32918 120000 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 179200 80928 180000 81048 6 io_in[2]
port 3 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 io_in[3]
port 4 nsew signal input
rlabel metal2 s 106278 119200 106334 120000 6 io_in[4]
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_in[5]
port 6 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 io_in[6]
port 7 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 io_in[7]
port 8 nsew signal input
rlabel metal2 s 142986 119200 143042 120000 6 io_out[0]
port 9 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 io_out[1]
port 10 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 io_out[2]
port 11 nsew signal output
rlabel metal2 s 179694 119200 179750 120000 6 io_out[3]
port 12 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 io_out[4]
port 13 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 io_out[5]
port 14 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[6]
port 15 nsew signal output
rlabel metal3 s 179200 3408 180000 3528 6 io_out[7]
port 16 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5360614
string GDS_FILE /home/runner/work/tiny_user_project/tiny_user_project/openlane/user_module/runs/22_09_06_09_12/results/signoff/user_module_334445762078310996.magic.gds
string GDS_START 23792
<< end >>

