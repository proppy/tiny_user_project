VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 170.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 9.560 150.000 10.160 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 111.560 150.000 112.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 121.760 150.000 122.360 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 131.960 150.000 132.560 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 142.160 150.000 142.760 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 152.360 150.000 152.960 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 166.000 146.650 170.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 166.000 130.090 170.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 166.000 113.530 170.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 166.000 96.970 170.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 166.000 80.410 170.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 19.760 150.000 20.360 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 166.000 63.850 170.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 166.000 47.290 170.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 166.000 30.730 170.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 166.000 14.170 170.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 29.960 150.000 30.560 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.160 150.000 40.760 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 50.360 150.000 50.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 60.560 150.000 61.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 70.760 150.000 71.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 80.960 150.000 81.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.160 150.000 91.760 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 101.360 150.000 101.960 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 16.360 150.000 16.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 118.360 150.000 118.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 128.560 150.000 129.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 138.760 150.000 139.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 148.960 150.000 149.560 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 159.160 150.000 159.760 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 166.000 135.610 170.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 166.000 119.050 170.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 166.000 102.490 170.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 166.000 85.930 170.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 166.000 69.370 170.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 26.560 150.000 27.160 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 166.000 52.810 170.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 166.000 36.250 170.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 166.000 19.690 170.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 166.000 3.130 170.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 36.760 150.000 37.360 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 46.960 150.000 47.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.160 150.000 57.760 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 67.360 150.000 67.960 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 77.560 150.000 78.160 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 87.760 150.000 88.360 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 97.960 150.000 98.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.160 150.000 108.760 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 12.960 150.000 13.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 114.960 150.000 115.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.160 150.000 125.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 135.360 150.000 135.960 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 145.560 150.000 146.160 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 155.760 150.000 156.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 166.000 141.130 170.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 166.000 124.570 170.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 166.000 108.010 170.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 166.000 91.450 170.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 166.000 74.890 170.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.160 150.000 23.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 166.000 58.330 170.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 166.000 41.770 170.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 166.000 25.210 170.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 166.000 8.650 170.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 33.360 150.000 33.960 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.560 150.000 44.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 53.760 150.000 54.360 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 63.960 150.000 64.560 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.160 150.000 74.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 84.360 150.000 84.960 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 94.560 150.000 95.160 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 104.760 150.000 105.360 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 158.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 158.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 158.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 157.845 ;
      LAYER met1 ;
        RECT 2.830 10.640 145.240 158.000 ;
      LAYER met2 ;
        RECT 3.410 165.720 8.090 166.000 ;
        RECT 8.930 165.720 13.610 166.000 ;
        RECT 14.450 165.720 19.130 166.000 ;
        RECT 19.970 165.720 24.650 166.000 ;
        RECT 25.490 165.720 30.170 166.000 ;
        RECT 31.010 165.720 35.690 166.000 ;
        RECT 36.530 165.720 41.210 166.000 ;
        RECT 42.050 165.720 46.730 166.000 ;
        RECT 47.570 165.720 52.250 166.000 ;
        RECT 53.090 165.720 57.770 166.000 ;
        RECT 58.610 165.720 63.290 166.000 ;
        RECT 64.130 165.720 68.810 166.000 ;
        RECT 69.650 165.720 74.330 166.000 ;
        RECT 75.170 165.720 79.850 166.000 ;
        RECT 80.690 165.720 85.370 166.000 ;
        RECT 86.210 165.720 90.890 166.000 ;
        RECT 91.730 165.720 96.410 166.000 ;
        RECT 97.250 165.720 101.930 166.000 ;
        RECT 102.770 165.720 107.450 166.000 ;
        RECT 108.290 165.720 112.970 166.000 ;
        RECT 113.810 165.720 118.490 166.000 ;
        RECT 119.330 165.720 124.010 166.000 ;
        RECT 124.850 165.720 129.530 166.000 ;
        RECT 130.370 165.720 135.050 166.000 ;
        RECT 135.890 165.720 140.570 166.000 ;
        RECT 141.410 165.720 145.210 166.000 ;
        RECT 2.860 10.695 145.210 165.720 ;
      LAYER met3 ;
        RECT 4.000 158.760 145.600 159.625 ;
        RECT 4.000 156.760 146.890 158.760 ;
        RECT 4.000 155.400 145.600 156.760 ;
        RECT 4.400 155.360 145.600 155.400 ;
        RECT 4.400 154.000 146.890 155.360 ;
        RECT 4.000 153.360 146.890 154.000 ;
        RECT 4.000 152.000 145.600 153.360 ;
        RECT 4.400 151.960 145.600 152.000 ;
        RECT 4.400 150.600 146.890 151.960 ;
        RECT 4.000 149.960 146.890 150.600 ;
        RECT 4.000 148.600 145.600 149.960 ;
        RECT 4.400 148.560 145.600 148.600 ;
        RECT 4.400 147.200 146.890 148.560 ;
        RECT 4.000 146.560 146.890 147.200 ;
        RECT 4.000 145.200 145.600 146.560 ;
        RECT 4.400 145.160 145.600 145.200 ;
        RECT 4.400 143.800 146.890 145.160 ;
        RECT 4.000 143.160 146.890 143.800 ;
        RECT 4.000 141.800 145.600 143.160 ;
        RECT 4.400 141.760 145.600 141.800 ;
        RECT 4.400 140.400 146.890 141.760 ;
        RECT 4.000 139.760 146.890 140.400 ;
        RECT 4.000 138.400 145.600 139.760 ;
        RECT 4.400 138.360 145.600 138.400 ;
        RECT 4.400 137.000 146.890 138.360 ;
        RECT 4.000 136.360 146.890 137.000 ;
        RECT 4.000 135.000 145.600 136.360 ;
        RECT 4.400 134.960 145.600 135.000 ;
        RECT 4.400 133.600 146.890 134.960 ;
        RECT 4.000 132.960 146.890 133.600 ;
        RECT 4.000 131.600 145.600 132.960 ;
        RECT 4.400 131.560 145.600 131.600 ;
        RECT 4.400 130.200 146.890 131.560 ;
        RECT 4.000 129.560 146.890 130.200 ;
        RECT 4.000 128.200 145.600 129.560 ;
        RECT 4.400 128.160 145.600 128.200 ;
        RECT 4.400 126.800 146.890 128.160 ;
        RECT 4.000 126.160 146.890 126.800 ;
        RECT 4.000 124.800 145.600 126.160 ;
        RECT 4.400 124.760 145.600 124.800 ;
        RECT 4.400 123.400 146.890 124.760 ;
        RECT 4.000 122.760 146.890 123.400 ;
        RECT 4.000 121.400 145.600 122.760 ;
        RECT 4.400 121.360 145.600 121.400 ;
        RECT 4.400 120.000 146.890 121.360 ;
        RECT 4.000 119.360 146.890 120.000 ;
        RECT 4.000 118.000 145.600 119.360 ;
        RECT 4.400 117.960 145.600 118.000 ;
        RECT 4.400 116.600 146.890 117.960 ;
        RECT 4.000 115.960 146.890 116.600 ;
        RECT 4.000 114.600 145.600 115.960 ;
        RECT 4.400 114.560 145.600 114.600 ;
        RECT 4.400 113.200 146.890 114.560 ;
        RECT 4.000 112.560 146.890 113.200 ;
        RECT 4.000 111.200 145.600 112.560 ;
        RECT 4.400 111.160 145.600 111.200 ;
        RECT 4.400 109.800 146.890 111.160 ;
        RECT 4.000 109.160 146.890 109.800 ;
        RECT 4.000 107.800 145.600 109.160 ;
        RECT 4.400 107.760 145.600 107.800 ;
        RECT 4.400 106.400 146.890 107.760 ;
        RECT 4.000 105.760 146.890 106.400 ;
        RECT 4.000 104.400 145.600 105.760 ;
        RECT 4.400 104.360 145.600 104.400 ;
        RECT 4.400 103.000 146.890 104.360 ;
        RECT 4.000 102.360 146.890 103.000 ;
        RECT 4.000 101.000 145.600 102.360 ;
        RECT 4.400 100.960 145.600 101.000 ;
        RECT 4.400 99.600 146.890 100.960 ;
        RECT 4.000 98.960 146.890 99.600 ;
        RECT 4.000 97.600 145.600 98.960 ;
        RECT 4.400 97.560 145.600 97.600 ;
        RECT 4.400 96.200 146.890 97.560 ;
        RECT 4.000 95.560 146.890 96.200 ;
        RECT 4.000 94.200 145.600 95.560 ;
        RECT 4.400 94.160 145.600 94.200 ;
        RECT 4.400 92.800 146.890 94.160 ;
        RECT 4.000 92.160 146.890 92.800 ;
        RECT 4.000 90.800 145.600 92.160 ;
        RECT 4.400 90.760 145.600 90.800 ;
        RECT 4.400 89.400 146.890 90.760 ;
        RECT 4.000 88.760 146.890 89.400 ;
        RECT 4.000 87.400 145.600 88.760 ;
        RECT 4.400 87.360 145.600 87.400 ;
        RECT 4.400 86.000 146.890 87.360 ;
        RECT 4.000 85.360 146.890 86.000 ;
        RECT 4.000 84.000 145.600 85.360 ;
        RECT 4.400 83.960 145.600 84.000 ;
        RECT 4.400 82.600 146.890 83.960 ;
        RECT 4.000 81.960 146.890 82.600 ;
        RECT 4.000 80.600 145.600 81.960 ;
        RECT 4.400 80.560 145.600 80.600 ;
        RECT 4.400 79.200 146.890 80.560 ;
        RECT 4.000 78.560 146.890 79.200 ;
        RECT 4.000 77.200 145.600 78.560 ;
        RECT 4.400 77.160 145.600 77.200 ;
        RECT 4.400 75.800 146.890 77.160 ;
        RECT 4.000 75.160 146.890 75.800 ;
        RECT 4.000 73.800 145.600 75.160 ;
        RECT 4.400 73.760 145.600 73.800 ;
        RECT 4.400 72.400 146.890 73.760 ;
        RECT 4.000 71.760 146.890 72.400 ;
        RECT 4.000 70.400 145.600 71.760 ;
        RECT 4.400 70.360 145.600 70.400 ;
        RECT 4.400 69.000 146.890 70.360 ;
        RECT 4.000 68.360 146.890 69.000 ;
        RECT 4.000 67.000 145.600 68.360 ;
        RECT 4.400 66.960 145.600 67.000 ;
        RECT 4.400 65.600 146.890 66.960 ;
        RECT 4.000 64.960 146.890 65.600 ;
        RECT 4.000 63.600 145.600 64.960 ;
        RECT 4.400 63.560 145.600 63.600 ;
        RECT 4.400 62.200 146.890 63.560 ;
        RECT 4.000 61.560 146.890 62.200 ;
        RECT 4.000 60.200 145.600 61.560 ;
        RECT 4.400 60.160 145.600 60.200 ;
        RECT 4.400 58.800 146.890 60.160 ;
        RECT 4.000 58.160 146.890 58.800 ;
        RECT 4.000 56.800 145.600 58.160 ;
        RECT 4.400 56.760 145.600 56.800 ;
        RECT 4.400 55.400 146.890 56.760 ;
        RECT 4.000 54.760 146.890 55.400 ;
        RECT 4.000 53.400 145.600 54.760 ;
        RECT 4.400 53.360 145.600 53.400 ;
        RECT 4.400 52.000 146.890 53.360 ;
        RECT 4.000 51.360 146.890 52.000 ;
        RECT 4.000 50.000 145.600 51.360 ;
        RECT 4.400 49.960 145.600 50.000 ;
        RECT 4.400 48.600 146.890 49.960 ;
        RECT 4.000 47.960 146.890 48.600 ;
        RECT 4.000 46.600 145.600 47.960 ;
        RECT 4.400 46.560 145.600 46.600 ;
        RECT 4.400 45.200 146.890 46.560 ;
        RECT 4.000 44.560 146.890 45.200 ;
        RECT 4.000 43.200 145.600 44.560 ;
        RECT 4.400 43.160 145.600 43.200 ;
        RECT 4.400 41.800 146.890 43.160 ;
        RECT 4.000 41.160 146.890 41.800 ;
        RECT 4.000 39.800 145.600 41.160 ;
        RECT 4.400 39.760 145.600 39.800 ;
        RECT 4.400 38.400 146.890 39.760 ;
        RECT 4.000 37.760 146.890 38.400 ;
        RECT 4.000 36.400 145.600 37.760 ;
        RECT 4.400 36.360 145.600 36.400 ;
        RECT 4.400 35.000 146.890 36.360 ;
        RECT 4.000 34.360 146.890 35.000 ;
        RECT 4.000 33.000 145.600 34.360 ;
        RECT 4.400 32.960 145.600 33.000 ;
        RECT 4.400 31.600 146.890 32.960 ;
        RECT 4.000 30.960 146.890 31.600 ;
        RECT 4.000 29.600 145.600 30.960 ;
        RECT 4.400 29.560 145.600 29.600 ;
        RECT 4.400 28.200 146.890 29.560 ;
        RECT 4.000 27.560 146.890 28.200 ;
        RECT 4.000 26.200 145.600 27.560 ;
        RECT 4.400 26.160 145.600 26.200 ;
        RECT 4.400 24.800 146.890 26.160 ;
        RECT 4.000 24.160 146.890 24.800 ;
        RECT 4.000 22.800 145.600 24.160 ;
        RECT 4.400 22.760 145.600 22.800 ;
        RECT 4.400 21.400 146.890 22.760 ;
        RECT 4.000 20.760 146.890 21.400 ;
        RECT 4.000 19.400 145.600 20.760 ;
        RECT 4.400 19.360 145.600 19.400 ;
        RECT 4.400 18.000 146.890 19.360 ;
        RECT 4.000 17.360 146.890 18.000 ;
        RECT 4.000 16.000 145.600 17.360 ;
        RECT 4.400 15.960 145.600 16.000 ;
        RECT 4.400 14.600 146.890 15.960 ;
        RECT 4.000 13.960 146.890 14.600 ;
        RECT 4.000 12.560 145.600 13.960 ;
        RECT 4.000 10.715 146.890 12.560 ;
  END
END tiny_user_project
END LIBRARY

