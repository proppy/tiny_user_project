magic
tech gf180mcuC
magscale 1 10
timestamp 1669350293
<< metal1 >>
rect 32274 46398 32286 46450
rect 32338 46447 32350 46450
rect 33170 46447 33182 46450
rect 32338 46401 33182 46447
rect 32338 46398 32350 46401
rect 33170 46398 33182 46401
rect 33234 46398 33246 46450
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 2270 45778 2322 45790
rect 2270 45714 2322 45726
rect 2942 45778 2994 45790
rect 2942 45714 2994 45726
rect 4286 45778 4338 45790
rect 4286 45714 4338 45726
rect 7646 45778 7698 45790
rect 7646 45714 7698 45726
rect 9662 45778 9714 45790
rect 9662 45714 9714 45726
rect 13582 45778 13634 45790
rect 13582 45714 13634 45726
rect 18398 45778 18450 45790
rect 18398 45714 18450 45726
rect 20414 45778 20466 45790
rect 20414 45714 20466 45726
rect 21758 45778 21810 45790
rect 21758 45714 21810 45726
rect 27134 45778 27186 45790
rect 27134 45714 27186 45726
rect 33182 45778 33234 45790
rect 33182 45714 33234 45726
rect 35870 45778 35922 45790
rect 35870 45714 35922 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 39902 45778 39954 45790
rect 39902 45714 39954 45726
rect 43262 45778 43314 45790
rect 43262 45714 43314 45726
rect 48078 45778 48130 45790
rect 48078 45714 48130 45726
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 1822 45330 1874 45342
rect 1822 45266 1874 45278
rect 2494 45330 2546 45342
rect 2494 45266 2546 45278
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 1822 44098 1874 44110
rect 1822 44034 1874 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 1822 42530 1874 42542
rect 1822 42466 1874 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 48078 40514 48130 40526
rect 48078 40450 48130 40462
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 1822 38946 1874 38958
rect 1822 38882 1874 38894
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 48078 37826 48130 37838
rect 48078 37762 48130 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 1822 37378 1874 37390
rect 1822 37314 1874 37326
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 48078 36258 48130 36270
rect 48078 36194 48130 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 1822 35810 1874 35822
rect 1822 35746 1874 35758
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 48078 34690 48130 34702
rect 48078 34626 48130 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 1822 33122 1874 33134
rect 1822 33058 1874 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 48078 32674 48130 32686
rect 48078 32610 48130 32622
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 48078 31554 48130 31566
rect 48078 31490 48130 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 48078 29538 48130 29550
rect 48078 29474 48130 29486
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 1822 28418 1874 28430
rect 1822 28354 1874 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 1822 26850 1874 26862
rect 1822 26786 1874 26798
rect 48078 26850 48130 26862
rect 48078 26786 48130 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 1822 24834 1874 24846
rect 1822 24770 1874 24782
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 48078 23714 48130 23726
rect 48078 23650 48130 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 1822 23266 1874 23278
rect 1822 23202 1874 23214
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 48078 22146 48130 22158
rect 48078 22082 48130 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 1822 19010 1874 19022
rect 1822 18946 1874 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 48078 18562 48130 18574
rect 48078 18498 48130 18510
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 1822 17554 1874 17566
rect 1822 17490 1874 17502
rect 48078 17442 48130 17454
rect 48078 17378 48130 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 1822 15874 1874 15886
rect 1822 15810 1874 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 1822 14306 1874 14318
rect 1822 14242 1874 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 48078 12850 48130 12862
rect 48078 12786 48130 12798
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 48078 12290 48130 12302
rect 48078 12226 48130 12238
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 1822 10722 1874 10734
rect 1822 10658 1874 10670
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 48078 9602 48130 9614
rect 48078 9538 48130 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 1822 9154 1874 9166
rect 1822 9090 1874 9102
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 48078 8034 48130 8046
rect 48078 7970 48130 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 1822 7586 1874 7598
rect 1822 7522 1874 7534
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 48078 6466 48130 6478
rect 48078 6402 48130 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 1822 4450 1874 4462
rect 1822 4386 1874 4398
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 1822 3330 1874 3342
rect 1822 3266 1874 3278
rect 2494 3330 2546 3342
rect 2494 3266 2546 3278
rect 3614 3330 3666 3342
rect 3614 3266 3666 3278
rect 5742 3330 5794 3342
rect 5742 3266 5794 3278
rect 9662 3330 9714 3342
rect 9662 3266 9714 3278
rect 14366 3330 14418 3342
rect 14366 3266 14418 3278
rect 15710 3330 15762 3342
rect 15710 3266 15762 3278
rect 17726 3330 17778 3342
rect 17726 3266 17778 3278
rect 21422 3330 21474 3342
rect 21422 3266 21474 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 29262 3330 29314 3342
rect 29262 3266 29314 3278
rect 31838 3330 31890 3342
rect 31838 3266 31890 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 41022 3330 41074 3342
rect 41022 3266 41074 3278
rect 42590 3330 42642 3342
rect 42590 3266 42642 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 45950 3330 46002 3342
rect 45950 3266 46002 3278
rect 47406 3330 47458 3342
rect 47406 3266 47458 3278
rect 48078 3330 48130 3342
rect 48078 3266 48130 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
rect 40338 1822 40350 1874
rect 40402 1871 40414 1874
rect 41010 1871 41022 1874
rect 40402 1825 41022 1871
rect 40402 1822 40414 1825
rect 41010 1822 41022 1825
rect 41074 1822 41086 1874
rect 8754 1710 8766 1762
rect 8818 1759 8830 1762
rect 9650 1759 9662 1762
rect 8818 1713 9662 1759
rect 8818 1710 8830 1713
rect 9650 1710 9662 1713
rect 9714 1710 9726 1762
rect 20850 1710 20862 1762
rect 20914 1759 20926 1762
rect 21410 1759 21422 1762
rect 20914 1713 21422 1759
rect 20914 1710 20926 1713
rect 21410 1710 21422 1713
rect 21474 1710 21486 1762
<< via1 >>
rect 32286 46398 32338 46450
rect 33182 46398 33234 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 2270 45726 2322 45778
rect 2942 45726 2994 45778
rect 4286 45726 4338 45778
rect 7646 45726 7698 45778
rect 9662 45726 9714 45778
rect 13582 45726 13634 45778
rect 18398 45726 18450 45778
rect 20414 45726 20466 45778
rect 21758 45726 21810 45778
rect 27134 45726 27186 45778
rect 33182 45726 33234 45778
rect 35870 45726 35922 45778
rect 37886 45726 37938 45778
rect 39902 45726 39954 45778
rect 43262 45726 43314 45778
rect 48078 45726 48130 45778
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 1822 45278 1874 45330
rect 2494 45278 2546 45330
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 1822 44046 1874 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 1822 42478 1874 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 48078 40462 48130 40514
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 1822 38894 1874 38946
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 48078 37774 48130 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 1822 37326 1874 37378
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 48078 36206 48130 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 1822 35758 1874 35810
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 48078 34638 48130 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 1822 33070 1874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 48078 32622 48130 32674
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 48078 31502 48130 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 1822 29934 1874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 48078 29486 48130 29538
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 1822 28366 1874 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1822 26798 1874 26850
rect 48078 26798 48130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 1822 24782 1874 24834
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 48078 23662 48130 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 1822 23214 1874 23266
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 48078 22094 48130 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 1822 21646 1874 21698
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 1822 18958 1874 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 48078 18510 48130 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 1822 17502 1874 17554
rect 48078 17390 48130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 1822 15822 1874 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14254 1874 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 48078 12798 48130 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 48078 12238 48130 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 1822 10670 1874 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 48078 9550 48130 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 1822 9102 1874 9154
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 48078 7982 48130 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 1822 7534 1874 7586
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 48078 6414 48130 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 1822 4398 1874 4450
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 1822 3278 1874 3330
rect 2494 3278 2546 3330
rect 3614 3278 3666 3330
rect 5742 3278 5794 3330
rect 9662 3278 9714 3330
rect 14366 3278 14418 3330
rect 15710 3278 15762 3330
rect 17726 3278 17778 3330
rect 21422 3278 21474 3330
rect 23102 3278 23154 3330
rect 26462 3278 26514 3330
rect 29262 3278 29314 3330
rect 31838 3278 31890 3330
rect 35198 3278 35250 3330
rect 38558 3278 38610 3330
rect 41022 3278 41074 3330
rect 42590 3278 42642 3330
rect 43934 3278 43986 3330
rect 45950 3278 46002 3330
rect 47406 3278 47458 3330
rect 48078 3278 48130 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 40350 1822 40402 1874
rect 41022 1822 41074 1874
rect 8766 1710 8818 1762
rect 9662 1710 9714 1762
rect 20862 1710 20914 1762
rect 21422 1710 21474 1762
<< metal2 >>
rect 672 49200 784 49800
rect 1036 49308 1876 49364
rect 700 49140 756 49200
rect 1036 49140 1092 49308
rect 700 49084 1092 49140
rect 1820 45330 1876 49308
rect 2016 49200 2128 49800
rect 4032 49200 4144 49800
rect 6048 49200 6160 49800
rect 7392 49200 7504 49800
rect 9408 49200 9520 49800
rect 11424 49200 11536 49800
rect 12768 49200 12880 49800
rect 14784 49200 14896 49800
rect 16128 49200 16240 49800
rect 18144 49200 18256 49800
rect 20160 49200 20272 49800
rect 21504 49200 21616 49800
rect 23520 49200 23632 49800
rect 25536 49200 25648 49800
rect 26880 49200 26992 49800
rect 28896 49200 29008 49800
rect 30912 49200 31024 49800
rect 32256 49200 32368 49800
rect 34272 49200 34384 49800
rect 35616 49200 35728 49800
rect 37632 49200 37744 49800
rect 39648 49200 39760 49800
rect 40992 49200 41104 49800
rect 43008 49200 43120 49800
rect 45024 49200 45136 49800
rect 46368 49200 46480 49800
rect 48384 49200 48496 49800
rect 49728 49200 49840 49800
rect 2044 45780 2100 49200
rect 3388 49140 3444 49150
rect 3388 47012 3444 49084
rect 2940 46956 3444 47012
rect 2268 45780 2324 45790
rect 2044 45778 2324 45780
rect 2044 45726 2270 45778
rect 2322 45726 2324 45778
rect 2044 45724 2324 45726
rect 2268 45714 2324 45724
rect 2492 45780 2548 45790
rect 1820 45278 1822 45330
rect 1874 45278 1876 45330
rect 1820 45266 1876 45278
rect 2492 45330 2548 45724
rect 2940 45778 2996 46956
rect 2940 45726 2942 45778
rect 2994 45726 2996 45778
rect 2940 45714 2996 45726
rect 4060 45780 4116 49200
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45780 4340 45790
rect 4060 45778 4340 45780
rect 4060 45726 4286 45778
rect 4338 45726 4340 45778
rect 4060 45724 4340 45726
rect 7420 45780 7476 49200
rect 7644 45780 7700 45790
rect 7420 45778 7700 45780
rect 7420 45726 7646 45778
rect 7698 45726 7700 45778
rect 7420 45724 7700 45726
rect 9436 45780 9492 49200
rect 9660 45780 9716 45790
rect 9436 45778 9716 45780
rect 9436 45726 9662 45778
rect 9714 45726 9716 45778
rect 9436 45724 9716 45726
rect 4284 45714 4340 45724
rect 7644 45714 7700 45724
rect 9660 45714 9716 45724
rect 12796 45780 12852 49200
rect 12796 45714 12852 45724
rect 13580 45780 13636 45790
rect 18172 45780 18228 49200
rect 18396 45780 18452 45790
rect 18172 45778 18452 45780
rect 18172 45726 18398 45778
rect 18450 45726 18452 45778
rect 18172 45724 18452 45726
rect 20188 45780 20244 49200
rect 20412 45780 20468 45790
rect 20188 45778 20468 45780
rect 20188 45726 20414 45778
rect 20466 45726 20468 45778
rect 20188 45724 20468 45726
rect 21532 45780 21588 49200
rect 21756 45780 21812 45790
rect 21532 45778 21812 45780
rect 21532 45726 21758 45778
rect 21810 45726 21812 45778
rect 21532 45724 21812 45726
rect 26908 45780 26964 49200
rect 32284 46450 32340 49200
rect 32284 46398 32286 46450
rect 32338 46398 32340 46450
rect 32284 46386 32340 46398
rect 33180 46450 33236 46462
rect 33180 46398 33182 46450
rect 33234 46398 33236 46450
rect 27132 45780 27188 45790
rect 26908 45778 27188 45780
rect 26908 45726 27134 45778
rect 27186 45726 27188 45778
rect 26908 45724 27188 45726
rect 13580 45686 13636 45724
rect 18396 45714 18452 45724
rect 20412 45714 20468 45724
rect 21756 45714 21812 45724
rect 27132 45714 27188 45724
rect 33180 45778 33236 46398
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 33180 45726 33182 45778
rect 33234 45726 33236 45778
rect 33180 45714 33236 45726
rect 35644 45780 35700 49200
rect 35868 45780 35924 45790
rect 35644 45778 35924 45780
rect 35644 45726 35870 45778
rect 35922 45726 35924 45778
rect 35644 45724 35924 45726
rect 37660 45780 37716 49200
rect 37884 45780 37940 45790
rect 37660 45778 37940 45780
rect 37660 45726 37886 45778
rect 37938 45726 37940 45778
rect 37660 45724 37940 45726
rect 39676 45780 39732 49200
rect 39900 45780 39956 45790
rect 39676 45778 39956 45780
rect 39676 45726 39902 45778
rect 39954 45726 39956 45778
rect 39676 45724 39956 45726
rect 43036 45780 43092 49200
rect 43260 45780 43316 45790
rect 43036 45778 43316 45780
rect 43036 45726 43262 45778
rect 43314 45726 43316 45778
rect 43036 45724 43316 45726
rect 35868 45714 35924 45724
rect 37884 45714 37940 45724
rect 39900 45714 39956 45724
rect 43260 45714 43316 45724
rect 48076 45780 48132 45790
rect 48412 45780 48468 49200
rect 48076 45778 48468 45780
rect 48076 45726 48078 45778
rect 48130 45726 48468 45778
rect 48076 45724 48468 45726
rect 48076 45714 48132 45724
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 2492 45278 2494 45330
rect 2546 45278 2548 45330
rect 2492 45266 2548 45278
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 1820 44098 1876 44110
rect 1820 44046 1822 44098
rect 1874 44046 1876 44098
rect 1820 43764 1876 44046
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 1820 43698 1876 43708
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 1820 42530 1876 42542
rect 1820 42478 1822 42530
rect 1874 42478 1876 42530
rect 1820 42420 1876 42478
rect 1820 42354 1876 42364
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 48076 40514 48132 40526
rect 48076 40462 48078 40514
rect 48130 40462 48132 40514
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 48076 39732 48132 40462
rect 48076 39666 48132 39676
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 1820 38946 1876 38958
rect 1820 38894 1822 38946
rect 1874 38894 1876 38946
rect 1820 38388 1876 38894
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 1820 38322 1876 38332
rect 48076 37826 48132 37838
rect 48076 37774 48078 37826
rect 48130 37774 48132 37826
rect 48076 37716 48132 37774
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 48076 37650 48132 37660
rect 19836 37594 20100 37604
rect 1820 37378 1876 37390
rect 1820 37326 1822 37378
rect 1874 37326 1876 37378
rect 1820 37044 1876 37326
rect 1820 36978 1876 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 48076 36258 48132 36270
rect 48076 36206 48078 36258
rect 48130 36206 48132 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 1820 35810 1876 35822
rect 1820 35758 1822 35810
rect 1874 35758 1876 35810
rect 1820 35028 1876 35758
rect 48076 35700 48132 36206
rect 48076 35634 48132 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 1820 34962 1876 34972
rect 48076 34690 48132 34702
rect 48076 34638 48078 34690
rect 48130 34638 48132 34690
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 48076 34356 48132 34638
rect 48076 34290 48132 34300
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 1820 33122 1876 33134
rect 1820 33070 1822 33122
rect 1874 33070 1876 33122
rect 1820 33012 1876 33070
rect 1820 32946 1876 32956
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 48076 32674 48132 32686
rect 48076 32622 48078 32674
rect 48130 32622 48132 32674
rect 48076 32340 48132 32622
rect 48076 32274 48132 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 48076 31554 48132 31566
rect 48076 31502 48078 31554
rect 48130 31502 48132 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 48076 30996 48132 31502
rect 48076 30930 48132 30940
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 1820 29986 1876 29998
rect 1820 29934 1822 29986
rect 1874 29934 1876 29986
rect 1820 29652 1876 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 1820 29586 1876 29596
rect 48076 29538 48132 29550
rect 48076 29486 48078 29538
rect 48130 29486 48132 29538
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 48076 28980 48132 29486
rect 48076 28914 48132 28924
rect 1820 28418 1876 28430
rect 1820 28366 1822 28418
rect 1874 28366 1876 28418
rect 1820 28308 1876 28366
rect 1820 28242 1876 28252
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 48076 26964 48132 26974
rect 1820 26850 1876 26862
rect 1820 26798 1822 26850
rect 1874 26798 1876 26850
rect 1820 26292 1876 26798
rect 48076 26850 48132 26908
rect 48076 26798 48078 26850
rect 48130 26798 48132 26850
rect 48076 26786 48132 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 1820 26226 1876 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 1820 24834 1876 24846
rect 1820 24782 1822 24834
rect 1874 24782 1876 24834
rect 1820 24276 1876 24782
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 1820 24210 1876 24220
rect 48076 23714 48132 23726
rect 48076 23662 48078 23714
rect 48130 23662 48132 23714
rect 48076 23604 48132 23662
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 48076 23538 48132 23548
rect 19836 23482 20100 23492
rect 1820 23266 1876 23278
rect 1820 23214 1822 23266
rect 1874 23214 1876 23266
rect 1820 22932 1876 23214
rect 1820 22866 1876 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 48076 22146 48132 22158
rect 48076 22094 48078 22146
rect 48130 22094 48132 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 1820 21698 1876 21710
rect 1820 21646 1822 21698
rect 1874 21646 1876 21698
rect 1820 20916 1876 21646
rect 48076 21588 48132 22094
rect 48076 21522 48132 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 1820 20850 1876 20860
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 1820 19010 1876 19022
rect 1820 18958 1822 19010
rect 1874 18958 1876 19010
rect 1820 18900 1876 18958
rect 1820 18834 1876 18844
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 48076 18562 48132 18574
rect 48076 18510 48078 18562
rect 48130 18510 48132 18562
rect 48076 18228 48132 18510
rect 48076 18162 48132 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 1820 17556 1876 17566
rect 1820 17462 1876 17500
rect 48076 17442 48132 17454
rect 48076 17390 48078 17442
rect 48130 17390 48132 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 48076 16884 48132 17390
rect 48076 16818 48132 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 1820 15874 1876 15886
rect 1820 15822 1822 15874
rect 1874 15822 1876 15874
rect 1820 15540 1876 15822
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 1820 15474 1876 15484
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 1820 14306 1876 14318
rect 1820 14254 1822 14306
rect 1874 14254 1876 14306
rect 1820 14196 1876 14254
rect 1820 14130 1876 14140
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 48076 12852 48132 12862
rect 48076 12758 48132 12796
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 48076 12290 48132 12302
rect 48076 12238 48078 12290
rect 48130 12238 48132 12290
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 48076 11508 48132 12238
rect 48076 11442 48132 11452
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 1820 10722 1876 10734
rect 1820 10670 1822 10722
rect 1874 10670 1876 10722
rect 1820 10164 1876 10670
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 1820 10098 1876 10108
rect 48076 9602 48132 9614
rect 48076 9550 48078 9602
rect 48130 9550 48132 9602
rect 48076 9492 48132 9550
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 48076 9426 48132 9436
rect 19836 9370 20100 9380
rect 1820 9154 1876 9166
rect 1820 9102 1822 9154
rect 1874 9102 1876 9154
rect 1820 8820 1876 9102
rect 1820 8754 1876 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 48076 8034 48132 8046
rect 48076 7982 48078 8034
rect 48130 7982 48132 8034
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 1820 7586 1876 7598
rect 1820 7534 1822 7586
rect 1874 7534 1876 7586
rect 1820 6804 1876 7534
rect 48076 7476 48132 7982
rect 48076 7410 48132 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 1820 6738 1876 6748
rect 48076 6466 48132 6478
rect 48076 6414 48078 6466
rect 48130 6414 48132 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 48076 6132 48132 6414
rect 48076 6066 48132 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 28 4452 84 4462
rect 28 800 84 4396
rect 1820 4452 1876 4462
rect 1820 4358 1876 4396
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 1820 3444 1876 3454
rect 1372 3332 1428 3342
rect 1372 800 1428 3276
rect 1820 3330 1876 3388
rect 1820 3278 1822 3330
rect 1874 3278 1876 3330
rect 1820 3266 1876 3278
rect 2492 3332 2548 3342
rect 3612 3332 3668 3342
rect 2492 3238 2548 3276
rect 3388 3330 3668 3332
rect 3388 3278 3614 3330
rect 3666 3278 3668 3330
rect 3388 3276 3668 3278
rect 3388 800 3444 3276
rect 3612 3266 3668 3276
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5740 3332 5796 3342
rect 5740 3238 5796 3276
rect 9660 3330 9716 3342
rect 14364 3332 14420 3342
rect 15708 3332 15764 3342
rect 17724 3332 17780 3342
rect 9660 3278 9662 3330
rect 9714 3278 9716 3330
rect 8764 1762 8820 1774
rect 8764 1710 8766 1762
rect 8818 1710 8820 1762
rect 8764 800 8820 1710
rect 9660 1762 9716 3278
rect 9660 1710 9662 1762
rect 9714 1710 9716 1762
rect 9660 1698 9716 1710
rect 14140 3330 14420 3332
rect 14140 3278 14366 3330
rect 14418 3278 14420 3330
rect 14140 3276 14420 3278
rect 14140 800 14196 3276
rect 14364 3266 14420 3276
rect 15484 3330 15764 3332
rect 15484 3278 15710 3330
rect 15762 3278 15764 3330
rect 15484 3276 15764 3278
rect 15484 800 15540 3276
rect 15708 3266 15764 3276
rect 17500 3330 17780 3332
rect 17500 3278 17726 3330
rect 17778 3278 17780 3330
rect 17500 3276 17780 3278
rect 17500 800 17556 3276
rect 17724 3266 17780 3276
rect 21420 3330 21476 3342
rect 23100 3332 23156 3342
rect 26460 3332 26516 3342
rect 21420 3278 21422 3330
rect 21474 3278 21476 3330
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 1762 20916 1774
rect 20860 1710 20862 1762
rect 20914 1710 20916 1762
rect 20860 800 20916 1710
rect 21420 1762 21476 3278
rect 21420 1710 21422 1762
rect 21474 1710 21476 1762
rect 21420 1698 21476 1710
rect 22876 3330 23156 3332
rect 22876 3278 23102 3330
rect 23154 3278 23156 3330
rect 22876 3276 23156 3278
rect 22876 800 22932 3276
rect 23100 3266 23156 3276
rect 26236 3330 26516 3332
rect 26236 3278 26462 3330
rect 26514 3278 26516 3330
rect 26236 3276 26516 3278
rect 26236 800 26292 3276
rect 26460 3266 26516 3276
rect 28252 3332 28308 3342
rect 28252 800 28308 3276
rect 29260 3332 29316 3342
rect 31836 3332 31892 3342
rect 35196 3332 35252 3342
rect 38556 3332 38612 3342
rect 29260 3238 29316 3276
rect 31612 3330 31892 3332
rect 31612 3278 31838 3330
rect 31890 3278 31892 3330
rect 31612 3276 31892 3278
rect 31612 800 31668 3276
rect 31836 3266 31892 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 41020 3330 41076 3342
rect 42588 3332 42644 3342
rect 43932 3332 43988 3342
rect 45948 3332 46004 3342
rect 41020 3278 41022 3330
rect 41074 3278 41076 3330
rect 40348 1874 40404 1886
rect 40348 1822 40350 1874
rect 40402 1822 40404 1874
rect 40348 800 40404 1822
rect 41020 1874 41076 3278
rect 41020 1822 41022 1874
rect 41074 1822 41076 1874
rect 41020 1810 41076 1822
rect 42364 3330 42644 3332
rect 42364 3278 42590 3330
rect 42642 3278 42644 3330
rect 42364 3276 42644 3278
rect 42364 800 42420 3276
rect 42588 3266 42644 3276
rect 43708 3330 43988 3332
rect 43708 3278 43934 3330
rect 43986 3278 43988 3330
rect 43708 3276 43988 3278
rect 43708 800 43764 3276
rect 43932 3266 43988 3276
rect 45724 3330 46004 3332
rect 45724 3278 45950 3330
rect 46002 3278 46004 3330
rect 45724 3276 46004 3278
rect 45724 800 45780 3276
rect 45948 3266 46004 3276
rect 47404 3330 47460 3342
rect 47404 3278 47406 3330
rect 47458 3278 47460 3330
rect 47404 2100 47460 3278
rect 47404 2034 47460 2044
rect 48076 3330 48132 3342
rect 48076 3278 48078 3330
rect 48130 3278 48132 3330
rect 0 200 112 800
rect 1344 200 1456 800
rect 3360 200 3472 800
rect 4704 200 4816 800
rect 6720 200 6832 800
rect 8736 200 8848 800
rect 10080 200 10192 800
rect 12096 200 12208 800
rect 14112 200 14224 800
rect 15456 200 15568 800
rect 17472 200 17584 800
rect 18816 200 18928 800
rect 20832 200 20944 800
rect 22848 200 22960 800
rect 24192 200 24304 800
rect 26208 200 26320 800
rect 28224 200 28336 800
rect 29568 200 29680 800
rect 31584 200 31696 800
rect 33600 200 33712 800
rect 34944 200 35056 800
rect 36960 200 37072 800
rect 38304 200 38416 800
rect 40320 200 40432 800
rect 42336 200 42448 800
rect 43680 200 43792 800
rect 45696 200 45808 800
rect 47712 200 47824 800
rect 48076 756 48132 3278
rect 48076 690 48132 700
rect 49056 200 49168 800
<< via2 >>
rect 3388 49084 3444 49140
rect 2492 45724 2548 45780
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 12796 45724 12852 45780
rect 13580 45778 13636 45780
rect 13580 45726 13582 45778
rect 13582 45726 13634 45778
rect 13634 45726 13636 45778
rect 13580 45724 13636 45726
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 1820 43708 1876 43764
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 1820 42364 1876 42420
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 48076 39676 48132 39732
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 1820 38332 1876 38388
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 48076 37660 48132 37716
rect 20044 37604 20100 37606
rect 1820 36988 1876 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 48076 35644 48132 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 1820 34972 1876 35028
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 48076 34300 48132 34356
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 1820 32956 1876 33012
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 48076 32284 48132 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 48076 30940 48132 30996
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 1820 29596 1876 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 48076 28924 48132 28980
rect 1820 28252 1876 28308
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 48076 26908 48132 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 1820 26236 1876 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 1820 24220 1876 24276
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 48076 23548 48132 23604
rect 20044 23492 20100 23494
rect 1820 22876 1876 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 48076 21532 48132 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 1820 20860 1876 20916
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 1820 18844 1876 18900
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 48076 18172 48132 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 1820 17554 1876 17556
rect 1820 17502 1822 17554
rect 1822 17502 1874 17554
rect 1874 17502 1876 17554
rect 1820 17500 1876 17502
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 48076 16828 48132 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 1820 15484 1876 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 1820 14140 1876 14196
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 48076 12850 48132 12852
rect 48076 12798 48078 12850
rect 48078 12798 48130 12850
rect 48130 12798 48132 12850
rect 48076 12796 48132 12798
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 48076 11452 48132 11508
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 1820 10108 1876 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 48076 9436 48132 9492
rect 20044 9380 20100 9382
rect 1820 8764 1876 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 48076 7420 48132 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 1820 6748 1876 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 48076 6076 48132 6132
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 28 4396 84 4452
rect 1820 4450 1876 4452
rect 1820 4398 1822 4450
rect 1822 4398 1874 4450
rect 1874 4398 1876 4450
rect 1820 4396 1876 4398
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 1820 3388 1876 3444
rect 1372 3276 1428 3332
rect 2492 3330 2548 3332
rect 2492 3278 2494 3330
rect 2494 3278 2546 3330
rect 2546 3278 2548 3330
rect 2492 3276 2548 3278
rect 4732 3276 4788 3332
rect 5740 3330 5796 3332
rect 5740 3278 5742 3330
rect 5742 3278 5794 3330
rect 5794 3278 5796 3330
rect 5740 3276 5796 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 28252 3276 28308 3332
rect 29260 3330 29316 3332
rect 29260 3278 29262 3330
rect 29262 3278 29314 3330
rect 29314 3278 29316 3330
rect 29260 3276 29316 3278
rect 47404 2044 47460 2100
rect 48076 700 48132 756
<< metal3 >>
rect 200 49140 800 49168
rect 200 49084 3388 49140
rect 3444 49084 3454 49140
rect 200 49056 800 49084
rect 49200 48384 49800 48496
rect 200 47712 800 47824
rect 49200 46368 49800 46480
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 200 45780 800 45808
rect 200 45724 2492 45780
rect 2548 45724 2558 45780
rect 12786 45724 12796 45780
rect 12852 45724 13580 45780
rect 13636 45724 13646 45780
rect 200 45696 800 45724
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 49200 45024 49800 45136
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 200 43764 800 43792
rect 200 43708 1820 43764
rect 1876 43708 1886 43764
rect 200 43680 800 43708
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 49200 43008 49800 43120
rect 200 42420 800 42448
rect 200 42364 1820 42420
rect 1876 42364 1886 42420
rect 200 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 49200 40992 49800 41104
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 200 40320 800 40432
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 49200 39732 49800 39760
rect 48066 39676 48076 39732
rect 48132 39676 49800 39732
rect 49200 39648 49800 39676
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 200 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 200 38332 1820 38388
rect 1876 38332 1886 38388
rect 200 38304 800 38332
rect 49200 37716 49800 37744
rect 48066 37660 48076 37716
rect 48132 37660 49800 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 49200 37632 49800 37660
rect 200 37044 800 37072
rect 200 36988 1820 37044
rect 1876 36988 1886 37044
rect 200 36960 800 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 49200 35700 49800 35728
rect 48066 35644 48076 35700
rect 48132 35644 49800 35700
rect 49200 35616 49800 35644
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 200 35028 800 35056
rect 200 34972 1820 35028
rect 1876 34972 1886 35028
rect 200 34944 800 34972
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 49200 34356 49800 34384
rect 48066 34300 48076 34356
rect 48132 34300 49800 34356
rect 49200 34272 49800 34300
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 200 33012 800 33040
rect 200 32956 1820 33012
rect 1876 32956 1886 33012
rect 200 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 49200 32340 49800 32368
rect 48066 32284 48076 32340
rect 48132 32284 49800 32340
rect 49200 32256 49800 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 200 31584 800 31696
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 49200 30996 49800 31024
rect 48066 30940 48076 30996
rect 48132 30940 49800 30996
rect 49200 30912 49800 30940
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 200 29652 800 29680
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 200 29568 800 29596
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 49200 28980 49800 29008
rect 48066 28924 48076 28980
rect 48132 28924 49800 28980
rect 49200 28896 49800 28924
rect 200 28308 800 28336
rect 200 28252 1820 28308
rect 1876 28252 1886 28308
rect 200 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 49200 26964 49800 26992
rect 48066 26908 48076 26964
rect 48132 26908 49800 26964
rect 49200 26880 49800 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 200 26292 800 26320
rect 200 26236 1820 26292
rect 1876 26236 1886 26292
rect 200 26208 800 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 49200 25536 49800 25648
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 200 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 200 24220 1820 24276
rect 1876 24220 1886 24276
rect 200 24192 800 24220
rect 49200 23604 49800 23632
rect 48066 23548 48076 23604
rect 48132 23548 49800 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 49200 23520 49800 23548
rect 200 22932 800 22960
rect 200 22876 1820 22932
rect 1876 22876 1886 22932
rect 200 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 49200 21588 49800 21616
rect 48066 21532 48076 21588
rect 48132 21532 49800 21588
rect 49200 21504 49800 21532
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 200 20916 800 20944
rect 200 20860 1820 20916
rect 1876 20860 1886 20916
rect 200 20832 800 20860
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 49200 20160 49800 20272
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 200 18900 800 18928
rect 200 18844 1820 18900
rect 1876 18844 1886 18900
rect 200 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 49200 18228 49800 18256
rect 48066 18172 48076 18228
rect 48132 18172 49800 18228
rect 49200 18144 49800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 200 17556 800 17584
rect 200 17500 1820 17556
rect 1876 17500 1886 17556
rect 200 17472 800 17500
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 49200 16884 49800 16912
rect 48066 16828 48076 16884
rect 48132 16828 49800 16884
rect 49200 16800 49800 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 200 15540 800 15568
rect 200 15484 1820 15540
rect 1876 15484 1886 15540
rect 200 15456 800 15484
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 49200 14784 49800 14896
rect 200 14196 800 14224
rect 200 14140 1820 14196
rect 1876 14140 1886 14196
rect 200 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 49200 12852 49800 12880
rect 48066 12796 48076 12852
rect 48132 12796 49800 12852
rect 49200 12768 49800 12796
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 200 12096 800 12208
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 49200 11508 49800 11536
rect 48066 11452 48076 11508
rect 48132 11452 49800 11508
rect 49200 11424 49800 11452
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 200 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 200 10108 1820 10164
rect 1876 10108 1886 10164
rect 200 10080 800 10108
rect 49200 9492 49800 9520
rect 48066 9436 48076 9492
rect 48132 9436 49800 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 49200 9408 49800 9436
rect 200 8820 800 8848
rect 200 8764 1820 8820
rect 1876 8764 1886 8820
rect 200 8736 800 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 49200 7476 49800 7504
rect 48066 7420 48076 7476
rect 48132 7420 49800 7476
rect 49200 7392 49800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 200 6804 800 6832
rect 200 6748 1820 6804
rect 1876 6748 1886 6804
rect 200 6720 800 6748
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 49200 6132 49800 6160
rect 48066 6076 48076 6132
rect 48132 6076 49800 6132
rect 49200 6048 49800 6076
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 200 4704 800 4816
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 18 4396 28 4452
rect 84 4396 1820 4452
rect 1876 4396 1886 4452
rect 49200 4032 49800 4144
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 200 3444 800 3472
rect 200 3388 1820 3444
rect 1876 3388 1886 3444
rect 200 3360 800 3388
rect 1362 3276 1372 3332
rect 1428 3276 2492 3332
rect 2548 3276 2558 3332
rect 4722 3276 4732 3332
rect 4788 3276 5740 3332
rect 5796 3276 5806 3332
rect 28242 3276 28252 3332
rect 28308 3276 29260 3332
rect 29316 3276 29326 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 49200 2100 49800 2128
rect 47394 2044 47404 2100
rect 47460 2044 49800 2100
rect 49200 2016 49800 2044
rect 200 1344 800 1456
rect 49200 756 49800 784
rect 48066 700 48076 756
rect 48132 700 49800 756
rect 49200 672 49800 700
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17
timestamp 1663859327
transform 1 0 3248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 3920 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31
timestamp 1663859327
transform 1 0 4816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1663859327
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 6048 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58
timestamp 1663859327
transform 1 0 7840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66
timestamp 1663859327
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1663859327
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77
timestamp 1663859327
transform 1 0 9968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93
timestamp 1663859327
transform 1 0 11760 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101
timestamp 1663859327
transform 1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1663859327
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119
timestamp 1663859327
transform 1 0 14672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_131
timestamp 1663859327
transform 1 0 16016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1663859327
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1663859327
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1663859327
transform 1 0 17472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_149
timestamp 1663859327
transform 1 0 18032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_165
timestamp 1663859327
transform 1 0 19824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1663859327
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1663859327
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182
timestamp 1663859327
transform 1 0 21728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1663859327
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192
timestamp 1663859327
transform 1 0 22848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_197
timestamp 1663859327
transform 1 0 23408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_205
timestamp 1663859327
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1663859327
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1663859327
transform 1 0 25088 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1663859327
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_222
timestamp 1663859327
transform 1 0 26208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_227
timestamp 1663859327
transform 1 0 26768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_243
timestamp 1663859327
transform 1 0 28560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1663859327
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_252
timestamp 1663859327
transform 1 0 29568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_268
timestamp 1663859327
transform 1 0 31360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_270
timestamp 1663859327
transform 1 0 31584 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_275
timestamp 1663859327
transform 1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1663859327
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_282
timestamp 1663859327
transform 1 0 32928 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1663859327
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_300
timestamp 1663859327
transform 1 0 34944 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_305
timestamp 1663859327
transform 1 0 35504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1663859327
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_317
timestamp 1663859327
transform 1 0 36848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_325
timestamp 1663859327
transform 1 0 37744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1663859327
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_335
timestamp 1663859327
transform 1 0 38864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_343
timestamp 1663859327
transform 1 0 39760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1663859327
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1663859327
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1663859327
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_357
timestamp 1663859327
transform 1 0 41328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_365
timestamp 1663859327
transform 1 0 42224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_371
timestamp 1663859327
transform 1 0 42896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_383
timestamp 1663859327
transform 1 0 44240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1663859327
transform 1 0 44688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_395
timestamp 1663859327
transform 1 0 45584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_401
timestamp 1663859327
transform 1 0 46256 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_413
timestamp 1663859327
transform 1 0 47600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1663859327
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1663859327
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_7 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2128 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1663859327
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1663859327
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1663859327
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1663859327
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1663859327
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1663859327
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1663859327
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1663859327
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1663859327
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1663859327
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1663859327
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1663859327
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 41328 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1663859327
transform 1 0 44912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_405
timestamp 1663859327
transform 1 0 46704 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_413
timestamp 1663859327
transform 1 0 47600 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1663859327
transform 1 0 48048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1663859327
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1663859327
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1663859327
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1663859327
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1663859327
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1663859327
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1663859327
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1663859327
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1663859327
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1663859327
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1663859327
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1663859327
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1663859327
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1663859327
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1663859327
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1663859327
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1663859327
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1663859327
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1663859327
transform 1 0 45248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1663859327
transform 1 0 47040 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_416
timestamp 1663859327
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1663859327
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1663859327
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1663859327
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1663859327
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1663859327
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1663859327
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1663859327
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1663859327
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1663859327
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1663859327
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1663859327
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1663859327
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1663859327
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1663859327
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1663859327
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_357
timestamp 1663859327
transform 1 0 41328 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1663859327
transform 1 0 44912 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1663859327
transform 1 0 46704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1663859327
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1663859327
transform 1 0 48048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1663859327
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1663859327
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1663859327
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1663859327
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1663859327
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1663859327
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1663859327
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1663859327
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1663859327
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1663859327
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1663859327
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1663859327
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1663859327
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1663859327
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1663859327
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1663859327
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1663859327
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1663859327
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1663859327
transform 1 0 45248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_408
timestamp 1663859327
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_412
timestamp 1663859327
transform 1 0 47488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_414
timestamp 1663859327
transform 1 0 47712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_419
timestamp 1663859327
transform 1 0 48272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1663859327
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_7
timestamp 1663859327
transform 1 0 2128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1663859327
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1663859327
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1663859327
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1663859327
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1663859327
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1663859327
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1663859327
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1663859327
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1663859327
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1663859327
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1663859327
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1663859327
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1663859327
transform 1 0 41328 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1663859327
transform 1 0 44912 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1663859327
transform 1 0 46704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1663859327
transform 1 0 47600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1663859327
transform 1 0 48048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1663859327
transform 1 0 48272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1663859327
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1663859327
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1663859327
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1663859327
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1663859327
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1663859327
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1663859327
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1663859327
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1663859327
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1663859327
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1663859327
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1663859327
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1663859327
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1663859327
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1663859327
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1663859327
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1663859327
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_392
timestamp 1663859327
transform 1 0 45248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_408
timestamp 1663859327
transform 1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_412
timestamp 1663859327
transform 1 0 47488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_414
timestamp 1663859327
transform 1 0 47712 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1663859327
transform 1 0 48272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1663859327
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_7
timestamp 1663859327
transform 1 0 2128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1663859327
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1663859327
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1663859327
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1663859327
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1663859327
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1663859327
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1663859327
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1663859327
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1663859327
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1663859327
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1663859327
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1663859327
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1663859327
transform 1 0 41328 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_389
timestamp 1663859327
transform 1 0 44912 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_405
timestamp 1663859327
transform 1 0 46704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_413
timestamp 1663859327
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1663859327
transform 1 0 48048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1663859327
transform 1 0 48272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1663859327
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1663859327
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1663859327
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1663859327
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1663859327
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1663859327
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1663859327
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1663859327
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1663859327
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1663859327
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1663859327
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1663859327
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1663859327
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1663859327
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1663859327
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1663859327
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1663859327
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1663859327
transform 1 0 45248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_408
timestamp 1663859327
transform 1 0 47040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_412
timestamp 1663859327
transform 1 0 47488 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_414
timestamp 1663859327
transform 1 0 47712 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_419
timestamp 1663859327
transform 1 0 48272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1663859327
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_7
timestamp 1663859327
transform 1 0 2128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1663859327
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1663859327
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1663859327
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1663859327
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1663859327
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1663859327
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1663859327
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1663859327
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1663859327
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1663859327
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1663859327
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1663859327
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_357
timestamp 1663859327
transform 1 0 41328 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_389
timestamp 1663859327
transform 1 0 44912 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1663859327
transform 1 0 46704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1663859327
transform 1 0 47600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1663859327
transform 1 0 48048 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1663859327
transform 1 0 48272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1663859327
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1663859327
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1663859327
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1663859327
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1663859327
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1663859327
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1663859327
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1663859327
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1663859327
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1663859327
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1663859327
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1663859327
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1663859327
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1663859327
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1663859327
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1663859327
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1663859327
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1663859327
transform 1 0 45248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1663859327
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1663859327
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1663859327
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1663859327
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1663859327
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1663859327
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1663859327
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1663859327
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1663859327
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1663859327
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1663859327
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1663859327
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1663859327
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1663859327
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1663859327
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1663859327
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1663859327
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_357
timestamp 1663859327
transform 1 0 41328 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1663859327
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1663859327
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_413
timestamp 1663859327
transform 1 0 47600 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1663859327
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1663859327
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1663859327
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1663859327
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1663859327
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1663859327
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1663859327
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1663859327
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1663859327
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1663859327
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1663859327
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1663859327
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1663859327
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1663859327
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1663859327
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1663859327
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1663859327
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1663859327
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_392
timestamp 1663859327
transform 1 0 45248 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_408
timestamp 1663859327
transform 1 0 47040 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_412
timestamp 1663859327
transform 1 0 47488 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_414
timestamp 1663859327
transform 1 0 47712 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1663859327
transform 1 0 48272 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1663859327
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1663859327
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1663859327
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1663859327
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1663859327
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1663859327
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1663859327
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1663859327
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1663859327
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1663859327
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1663859327
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1663859327
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1663859327
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1663859327
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1663859327
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1663859327
transform 1 0 41328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_389
timestamp 1663859327
transform 1 0 44912 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_405
timestamp 1663859327
transform 1 0 46704 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1663859327
transform 1 0 47600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1663859327
transform 1 0 48048 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1663859327
transform 1 0 48272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1663859327
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_7
timestamp 1663859327
transform 1 0 2128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_23
timestamp 1663859327
transform 1 0 3920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1663859327
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1663859327
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1663859327
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1663859327
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1663859327
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1663859327
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1663859327
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1663859327
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1663859327
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1663859327
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1663859327
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1663859327
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1663859327
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1663859327
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1663859327
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1663859327
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_392
timestamp 1663859327
transform 1 0 45248 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1663859327
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1663859327
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1663859327
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1663859327
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1663859327
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1663859327
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1663859327
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1663859327
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1663859327
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1663859327
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1663859327
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1663859327
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1663859327
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1663859327
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1663859327
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1663859327
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1663859327
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_357
timestamp 1663859327
transform 1 0 41328 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_389
timestamp 1663859327
transform 1 0 44912 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_405
timestamp 1663859327
transform 1 0 46704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1663859327
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_417
timestamp 1663859327
transform 1 0 48048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1663859327
transform 1 0 48272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1663859327
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_7
timestamp 1663859327
transform 1 0 2128 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_23
timestamp 1663859327
transform 1 0 3920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_31
timestamp 1663859327
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1663859327
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1663859327
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1663859327
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1663859327
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1663859327
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1663859327
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1663859327
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1663859327
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1663859327
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1663859327
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1663859327
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1663859327
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1663859327
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1663859327
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1663859327
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_392
timestamp 1663859327
transform 1 0 45248 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1663859327
transform 1 0 47040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1663859327
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1663859327
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1663859327
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1663859327
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1663859327
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1663859327
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1663859327
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1663859327
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1663859327
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1663859327
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1663859327
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1663859327
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1663859327
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1663859327
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1663859327
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1663859327
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_357
timestamp 1663859327
transform 1 0 41328 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_389
timestamp 1663859327
transform 1 0 44912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_405
timestamp 1663859327
transform 1 0 46704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_413
timestamp 1663859327
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_417
timestamp 1663859327
transform 1 0 48048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1663859327
transform 1 0 48272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1663859327
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_7
timestamp 1663859327
transform 1 0 2128 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_23
timestamp 1663859327
transform 1 0 3920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_31
timestamp 1663859327
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1663859327
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1663859327
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1663859327
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1663859327
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1663859327
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1663859327
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1663859327
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1663859327
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1663859327
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1663859327
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1663859327
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1663859327
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1663859327
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1663859327
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1663859327
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_392
timestamp 1663859327
transform 1 0 45248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_408
timestamp 1663859327
transform 1 0 47040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_412
timestamp 1663859327
transform 1 0 47488 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_414
timestamp 1663859327
transform 1 0 47712 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_419
timestamp 1663859327
transform 1 0 48272 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1663859327
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1663859327
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1663859327
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1663859327
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1663859327
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1663859327
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1663859327
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1663859327
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1663859327
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1663859327
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1663859327
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1663859327
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1663859327
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1663859327
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1663859327
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_357
timestamp 1663859327
transform 1 0 41328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_389
timestamp 1663859327
transform 1 0 44912 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_405
timestamp 1663859327
transform 1 0 46704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_413
timestamp 1663859327
transform 1 0 47600 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1663859327
transform 1 0 48272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1663859327
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_7
timestamp 1663859327
transform 1 0 2128 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_23
timestamp 1663859327
transform 1 0 3920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_31
timestamp 1663859327
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1663859327
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1663859327
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1663859327
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1663859327
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1663859327
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1663859327
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1663859327
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1663859327
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1663859327
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1663859327
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1663859327
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1663859327
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1663859327
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1663859327
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1663859327
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_392
timestamp 1663859327
transform 1 0 45248 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_408
timestamp 1663859327
transform 1 0 47040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_416
timestamp 1663859327
transform 1 0 47936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1663859327
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1663859327
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1663859327
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1663859327
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1663859327
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1663859327
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1663859327
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1663859327
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1663859327
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1663859327
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1663859327
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1663859327
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1663859327
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1663859327
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1663859327
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1663859327
transform 1 0 41328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_389
timestamp 1663859327
transform 1 0 44912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_405
timestamp 1663859327
transform 1 0 46704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_413
timestamp 1663859327
transform 1 0 47600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_417
timestamp 1663859327
transform 1 0 48048 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1663859327
transform 1 0 48272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1663859327
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1663859327
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1663859327
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1663859327
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1663859327
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1663859327
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1663859327
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1663859327
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1663859327
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1663859327
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1663859327
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1663859327
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1663859327
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1663859327
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1663859327
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1663859327
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1663859327
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_392
timestamp 1663859327
transform 1 0 45248 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_408
timestamp 1663859327
transform 1 0 47040 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_416
timestamp 1663859327
transform 1 0 47936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1663859327
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_7
timestamp 1663859327
transform 1 0 2128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1663859327
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1663859327
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1663859327
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1663859327
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1663859327
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1663859327
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1663859327
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1663859327
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1663859327
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1663859327
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1663859327
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1663859327
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_357
timestamp 1663859327
transform 1 0 41328 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_389
timestamp 1663859327
transform 1 0 44912 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_405
timestamp 1663859327
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_413
timestamp 1663859327
transform 1 0 47600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_417
timestamp 1663859327
transform 1 0 48048 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1663859327
transform 1 0 48272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1663859327
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1663859327
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1663859327
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1663859327
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1663859327
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1663859327
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1663859327
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1663859327
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1663859327
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1663859327
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1663859327
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1663859327
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1663859327
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1663859327
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1663859327
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1663859327
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1663859327
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_392
timestamp 1663859327
transform 1 0 45248 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_408
timestamp 1663859327
transform 1 0 47040 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_412
timestamp 1663859327
transform 1 0 47488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_414
timestamp 1663859327
transform 1 0 47712 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1663859327
transform 1 0 48272 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1663859327
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_7
timestamp 1663859327
transform 1 0 2128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1663859327
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1663859327
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1663859327
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1663859327
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1663859327
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1663859327
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1663859327
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1663859327
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1663859327
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1663859327
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1663859327
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1663859327
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1663859327
transform 1 0 41328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_389
timestamp 1663859327
transform 1 0 44912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_405
timestamp 1663859327
transform 1 0 46704 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_413
timestamp 1663859327
transform 1 0 47600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1663859327
transform 1 0 48048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1663859327
transform 1 0 48272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1663859327
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1663859327
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1663859327
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1663859327
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1663859327
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1663859327
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1663859327
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1663859327
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1663859327
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1663859327
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1663859327
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1663859327
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1663859327
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1663859327
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1663859327
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1663859327
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1663859327
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_392
timestamp 1663859327
transform 1 0 45248 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_408
timestamp 1663859327
transform 1 0 47040 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_412
timestamp 1663859327
transform 1 0 47488 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_414
timestamp 1663859327
transform 1 0 47712 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1663859327
transform 1 0 48272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1663859327
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_7
timestamp 1663859327
transform 1 0 2128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1663859327
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1663859327
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1663859327
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1663859327
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1663859327
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1663859327
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1663859327
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1663859327
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1663859327
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1663859327
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1663859327
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1663859327
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1663859327
transform 1 0 41328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_389
timestamp 1663859327
transform 1 0 44912 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_405
timestamp 1663859327
transform 1 0 46704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1663859327
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1663859327
transform 1 0 48048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1663859327
transform 1 0 48272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1663859327
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1663859327
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1663859327
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1663859327
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1663859327
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1663859327
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1663859327
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1663859327
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1663859327
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1663859327
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1663859327
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1663859327
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1663859327
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1663859327
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1663859327
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1663859327
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1663859327
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_392
timestamp 1663859327
transform 1 0 45248 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_408
timestamp 1663859327
transform 1 0 47040 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_416
timestamp 1663859327
transform 1 0 47936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1663859327
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1663859327
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1663859327
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1663859327
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1663859327
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1663859327
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1663859327
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1663859327
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1663859327
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1663859327
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1663859327
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1663859327
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1663859327
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1663859327
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1663859327
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_357
timestamp 1663859327
transform 1 0 41328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_389
timestamp 1663859327
transform 1 0 44912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_405
timestamp 1663859327
transform 1 0 46704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_413
timestamp 1663859327
transform 1 0 47600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1663859327
transform 1 0 48048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1663859327
transform 1 0 48272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1663859327
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_7
timestamp 1663859327
transform 1 0 2128 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_23
timestamp 1663859327
transform 1 0 3920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_31
timestamp 1663859327
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1663859327
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1663859327
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1663859327
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1663859327
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1663859327
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1663859327
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1663859327
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1663859327
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1663859327
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1663859327
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1663859327
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1663859327
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1663859327
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1663859327
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1663859327
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_392
timestamp 1663859327
transform 1 0 45248 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_408
timestamp 1663859327
transform 1 0 47040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_412
timestamp 1663859327
transform 1 0 47488 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_414
timestamp 1663859327
transform 1 0 47712 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_419
timestamp 1663859327
transform 1 0 48272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1663859327
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1663859327
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1663859327
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1663859327
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1663859327
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1663859327
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1663859327
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1663859327
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1663859327
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1663859327
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1663859327
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1663859327
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1663859327
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1663859327
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1663859327
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_357
timestamp 1663859327
transform 1 0 41328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_389
timestamp 1663859327
transform 1 0 44912 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_405
timestamp 1663859327
transform 1 0 46704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_413
timestamp 1663859327
transform 1 0 47600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_417
timestamp 1663859327
transform 1 0 48048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1663859327
transform 1 0 48272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1663859327
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_7
timestamp 1663859327
transform 1 0 2128 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_23
timestamp 1663859327
transform 1 0 3920 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_31
timestamp 1663859327
transform 1 0 4816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1663859327
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1663859327
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1663859327
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1663859327
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1663859327
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1663859327
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1663859327
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1663859327
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1663859327
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1663859327
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1663859327
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1663859327
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1663859327
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1663859327
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1663859327
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_392
timestamp 1663859327
transform 1 0 45248 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_408
timestamp 1663859327
transform 1 0 47040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_416
timestamp 1663859327
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1663859327
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1663859327
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1663859327
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1663859327
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1663859327
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1663859327
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1663859327
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1663859327
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1663859327
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1663859327
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1663859327
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1663859327
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1663859327
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1663859327
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1663859327
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1663859327
transform 1 0 41328 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_389
timestamp 1663859327
transform 1 0 44912 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_405
timestamp 1663859327
transform 1 0 46704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_413
timestamp 1663859327
transform 1 0 47600 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1663859327
transform 1 0 48272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1663859327
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_7
timestamp 1663859327
transform 1 0 2128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_23
timestamp 1663859327
transform 1 0 3920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_31
timestamp 1663859327
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1663859327
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1663859327
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1663859327
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1663859327
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1663859327
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1663859327
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1663859327
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1663859327
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1663859327
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1663859327
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1663859327
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1663859327
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1663859327
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1663859327
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1663859327
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_392
timestamp 1663859327
transform 1 0 45248 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_408
timestamp 1663859327
transform 1 0 47040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_416
timestamp 1663859327
transform 1 0 47936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1663859327
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1663859327
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1663859327
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1663859327
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1663859327
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1663859327
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1663859327
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1663859327
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1663859327
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1663859327
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1663859327
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1663859327
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1663859327
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1663859327
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1663859327
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_357
timestamp 1663859327
transform 1 0 41328 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_389
timestamp 1663859327
transform 1 0 44912 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_405
timestamp 1663859327
transform 1 0 46704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_413
timestamp 1663859327
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_417
timestamp 1663859327
transform 1 0 48048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_419
timestamp 1663859327
transform 1 0 48272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1663859327
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1663859327
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1663859327
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1663859327
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1663859327
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1663859327
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1663859327
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1663859327
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1663859327
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1663859327
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1663859327
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1663859327
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1663859327
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1663859327
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1663859327
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1663859327
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1663859327
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_392
timestamp 1663859327
transform 1 0 45248 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_408
timestamp 1663859327
transform 1 0 47040 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_412
timestamp 1663859327
transform 1 0 47488 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_414
timestamp 1663859327
transform 1 0 47712 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_419
timestamp 1663859327
transform 1 0 48272 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1663859327
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1663859327
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1663859327
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1663859327
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1663859327
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1663859327
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1663859327
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1663859327
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1663859327
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1663859327
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1663859327
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1663859327
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1663859327
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1663859327
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1663859327
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_357
timestamp 1663859327
transform 1 0 41328 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_389
timestamp 1663859327
transform 1 0 44912 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_405
timestamp 1663859327
transform 1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_413
timestamp 1663859327
transform 1 0 47600 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1663859327
transform 1 0 48272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1663859327
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_7
timestamp 1663859327
transform 1 0 2128 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_23
timestamp 1663859327
transform 1 0 3920 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_31
timestamp 1663859327
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1663859327
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1663859327
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1663859327
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1663859327
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1663859327
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1663859327
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1663859327
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1663859327
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1663859327
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1663859327
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1663859327
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1663859327
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1663859327
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1663859327
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1663859327
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_392
timestamp 1663859327
transform 1 0 45248 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_408
timestamp 1663859327
transform 1 0 47040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_416
timestamp 1663859327
transform 1 0 47936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1663859327
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1663859327
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1663859327
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1663859327
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1663859327
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1663859327
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1663859327
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1663859327
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1663859327
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1663859327
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1663859327
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1663859327
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1663859327
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1663859327
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1663859327
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1663859327
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_389
timestamp 1663859327
transform 1 0 44912 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_405
timestamp 1663859327
transform 1 0 46704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_413
timestamp 1663859327
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_417
timestamp 1663859327
transform 1 0 48048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1663859327
transform 1 0 48272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1663859327
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1663859327
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1663859327
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1663859327
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1663859327
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1663859327
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1663859327
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1663859327
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1663859327
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1663859327
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1663859327
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1663859327
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1663859327
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1663859327
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1663859327
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1663859327
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1663859327
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_392
timestamp 1663859327
transform 1 0 45248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_408
timestamp 1663859327
transform 1 0 47040 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_412
timestamp 1663859327
transform 1 0 47488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_414
timestamp 1663859327
transform 1 0 47712 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_419
timestamp 1663859327
transform 1 0 48272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1663859327
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_7
timestamp 1663859327
transform 1 0 2128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1663859327
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1663859327
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1663859327
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1663859327
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1663859327
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1663859327
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1663859327
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1663859327
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1663859327
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1663859327
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1663859327
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1663859327
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_357
timestamp 1663859327
transform 1 0 41328 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_389
timestamp 1663859327
transform 1 0 44912 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_405
timestamp 1663859327
transform 1 0 46704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_413
timestamp 1663859327
transform 1 0 47600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_417
timestamp 1663859327
transform 1 0 48048 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1663859327
transform 1 0 48272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1663859327
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1663859327
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1663859327
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1663859327
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1663859327
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1663859327
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1663859327
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1663859327
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1663859327
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1663859327
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1663859327
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1663859327
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1663859327
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1663859327
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1663859327
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1663859327
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1663859327
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1663859327
transform 1 0 45248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_408
timestamp 1663859327
transform 1 0 47040 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_412
timestamp 1663859327
transform 1 0 47488 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_414
timestamp 1663859327
transform 1 0 47712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1663859327
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1663859327
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_7
timestamp 1663859327
transform 1 0 2128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1663859327
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1663859327
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1663859327
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1663859327
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1663859327
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1663859327
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1663859327
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1663859327
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1663859327
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1663859327
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1663859327
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1663859327
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_357
timestamp 1663859327
transform 1 0 41328 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_389
timestamp 1663859327
transform 1 0 44912 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_405
timestamp 1663859327
transform 1 0 46704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_413
timestamp 1663859327
transform 1 0 47600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_417
timestamp 1663859327
transform 1 0 48048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_419
timestamp 1663859327
transform 1 0 48272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1663859327
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1663859327
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1663859327
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1663859327
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1663859327
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1663859327
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1663859327
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1663859327
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1663859327
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1663859327
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1663859327
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1663859327
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1663859327
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1663859327
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1663859327
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1663859327
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1663859327
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1663859327
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_408
timestamp 1663859327
transform 1 0 47040 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_412
timestamp 1663859327
transform 1 0 47488 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_414
timestamp 1663859327
transform 1 0 47712 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_419
timestamp 1663859327
transform 1 0 48272 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1663859327
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_7
timestamp 1663859327
transform 1 0 2128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1663859327
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1663859327
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1663859327
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1663859327
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1663859327
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1663859327
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1663859327
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1663859327
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1663859327
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1663859327
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1663859327
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1663859327
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_357
timestamp 1663859327
transform 1 0 41328 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_389
timestamp 1663859327
transform 1 0 44912 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_405
timestamp 1663859327
transform 1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_413
timestamp 1663859327
transform 1 0 47600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_417
timestamp 1663859327
transform 1 0 48048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1663859327
transform 1 0 48272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1663859327
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1663859327
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1663859327
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1663859327
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1663859327
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1663859327
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1663859327
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1663859327
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1663859327
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1663859327
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1663859327
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1663859327
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1663859327
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1663859327
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1663859327
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1663859327
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1663859327
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1663859327
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_408
timestamp 1663859327
transform 1 0 47040 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_416
timestamp 1663859327
transform 1 0 47936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1663859327
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1663859327
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1663859327
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1663859327
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1663859327
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1663859327
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1663859327
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1663859327
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1663859327
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1663859327
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1663859327
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1663859327
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1663859327
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1663859327
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1663859327
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1663859327
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1663859327
transform 1 0 44912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1663859327
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_413
timestamp 1663859327
transform 1 0 47600 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1663859327
transform 1 0 48272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1663859327
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1663859327
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1663859327
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1663859327
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1663859327
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1663859327
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1663859327
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1663859327
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1663859327
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1663859327
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1663859327
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1663859327
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1663859327
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1663859327
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1663859327
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1663859327
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1663859327
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1663859327
transform 1 0 45248 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_408
timestamp 1663859327
transform 1 0 47040 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_416
timestamp 1663859327
transform 1 0 47936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1663859327
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1663859327
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1663859327
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1663859327
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1663859327
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1663859327
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1663859327
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1663859327
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1663859327
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1663859327
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1663859327
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1663859327
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1663859327
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1663859327
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1663859327
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1663859327
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1663859327
transform 1 0 44912 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1663859327
transform 1 0 46704 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1663859327
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1663859327
transform 1 0 48048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1663859327
transform 1 0 48272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1663859327
transform 1 0 1568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_7
timestamp 1663859327
transform 1 0 2128 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_23
timestamp 1663859327
transform 1 0 3920 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_31
timestamp 1663859327
transform 1 0 4816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1663859327
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1663859327
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1663859327
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1663859327
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1663859327
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1663859327
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1663859327
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1663859327
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1663859327
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1663859327
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1663859327
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1663859327
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1663859327
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1663859327
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1663859327
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1663859327
transform 1 0 45248 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_408
timestamp 1663859327
transform 1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_416
timestamp 1663859327
transform 1 0 47936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1663859327
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1663859327
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1663859327
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1663859327
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1663859327
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1663859327
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1663859327
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1663859327
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1663859327
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1663859327
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1663859327
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1663859327
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1663859327
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1663859327
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1663859327
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1663859327
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1663859327
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1663859327
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1663859327
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1663859327
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1663859327
transform 1 0 48272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1663859327
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_7
timestamp 1663859327
transform 1 0 2128 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_23
timestamp 1663859327
transform 1 0 3920 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_31
timestamp 1663859327
transform 1 0 4816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1663859327
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1663859327
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1663859327
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1663859327
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1663859327
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1663859327
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1663859327
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1663859327
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1663859327
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1663859327
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1663859327
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1663859327
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1663859327
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1663859327
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1663859327
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1663859327
transform 1 0 45248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1663859327
transform 1 0 47040 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_416
timestamp 1663859327
transform 1 0 47936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1663859327
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_7
timestamp 1663859327
transform 1 0 2128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_13
timestamp 1663859327
transform 1 0 2800 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_45
timestamp 1663859327
transform 1 0 6384 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_61
timestamp 1663859327
transform 1 0 8176 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1663859327
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1663859327
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1663859327
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1663859327
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1663859327
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1663859327
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1663859327
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1663859327
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1663859327
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1663859327
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1663859327
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1663859327
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1663859327
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1663859327
transform 1 0 41328 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_389
timestamp 1663859327
transform 1 0 44912 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_405
timestamp 1663859327
transform 1 0 46704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_413
timestamp 1663859327
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_417
timestamp 1663859327
transform 1 0 48048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1663859327
transform 1 0 48272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_2
timestamp 1663859327
transform 1 0 1568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_6
timestamp 1663859327
transform 1 0 2016 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_11
timestamp 1663859327
transform 1 0 2576 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_17
timestamp 1663859327
transform 1 0 3248 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1663859327
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1663859327
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_37
timestamp 1663859327
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_53
timestamp 1663859327
transform 1 0 7280 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_59
timestamp 1663859327
transform 1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_67
timestamp 1663859327
transform 1 0 8848 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1663859327
transform 1 0 9072 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_72
timestamp 1663859327
transform 1 0 9408 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_77
timestamp 1663859327
transform 1 0 9968 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_93
timestamp 1663859327
transform 1 0 11760 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1663859327
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_107
timestamp 1663859327
transform 1 0 13328 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_112
timestamp 1663859327
transform 1 0 13888 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_128
timestamp 1663859327
transform 1 0 15680 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_136
timestamp 1663859327
transform 1 0 16576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_142
timestamp 1663859327
transform 1 0 17248 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_150
timestamp 1663859327
transform 1 0 18144 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_155
timestamp 1663859327
transform 1 0 18704 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_163
timestamp 1663859327
transform 1 0 19600 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_167
timestamp 1663859327
transform 1 0 20048 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_173
timestamp 1663859327
transform 1 0 20720 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_177
timestamp 1663859327
transform 1 0 21168 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_185
timestamp 1663859327
transform 1 0 22064 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_201
timestamp 1663859327
transform 1 0 23856 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_209
timestamp 1663859327
transform 1 0 24752 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_212
timestamp 1663859327
transform 1 0 25088 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_228
timestamp 1663859327
transform 1 0 26880 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_233
timestamp 1663859327
transform 1 0 27440 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_241
timestamp 1663859327
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_247
timestamp 1663859327
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1663859327
transform 1 0 32592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_282
timestamp 1663859327
transform 1 0 32928 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_287
timestamp 1663859327
transform 1 0 33488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_303
timestamp 1663859327
transform 1 0 35280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_311
timestamp 1663859327
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_317
timestamp 1663859327
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_329
timestamp 1663859327
transform 1 0 38192 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_337
timestamp 1663859327
transform 1 0 39088 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_341
timestamp 1663859327
transform 1 0 39536 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_347
timestamp 1663859327
transform 1 0 40208 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1663859327
transform 1 0 40432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_352
timestamp 1663859327
transform 1 0 40768 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_368
timestamp 1663859327
transform 1 0 42560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_372
timestamp 1663859327
transform 1 0 43008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_377
timestamp 1663859327
transform 1 0 43568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_387
timestamp 1663859327
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_403
timestamp 1663859327
transform 1 0 46480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_411
timestamp 1663859327
transform 1 0 47376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1663859327
transform 1 0 48272 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1663859327
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1663859327
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1663859327
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1663859327
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1663859327
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1663859327
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1663859327
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1663859327
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1663859327
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1663859327
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1663859327
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1663859327
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1663859327
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1663859327
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1663859327
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1663859327
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1663859327
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1663859327
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1663859327
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1663859327
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1663859327
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1663859327
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1663859327
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1663859327
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1663859327
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1663859327
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1663859327
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1663859327
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1663859327
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1663859327
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1663859327
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1663859327
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1663859327
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1663859327
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1663859327
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1663859327
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1663859327
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1663859327
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1663859327
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1663859327
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1663859327
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1663859327
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1663859327
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1663859327
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1663859327
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1663859327
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1663859327
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1663859327
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1663859327
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1663859327
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1663859327
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1663859327
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1663859327
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1663859327
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1663859327
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1663859327
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1663859327
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1663859327
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1663859327
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1663859327
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1663859327
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1663859327
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1663859327
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1663859327
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1663859327
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1663859327
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1663859327
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1663859327
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1663859327
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1663859327
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1663859327
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1663859327
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1663859327
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1663859327
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1663859327
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1663859327
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1663859327
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1663859327
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1663859327
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1663859327
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1663859327
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1663859327
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1663859327
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1663859327
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1663859327
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1663859327
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1663859327
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1663859327
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1663859327
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1663859327
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1663859327
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1663859327
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1663859327
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1663859327
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1663859327
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1663859327
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1663859327
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1663859327
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1663859327
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1663859327
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1663859327
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1663859327
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1663859327
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1663859327
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1663859327
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1663859327
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1663859327
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1663859327
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1663859327
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1663859327
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1663859327
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1663859327
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1663859327
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1663859327
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1663859327
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1663859327
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1663859327
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1663859327
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1663859327
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1663859327
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1663859327
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1663859327
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1663859327
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1663859327
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1663859327
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1663859327
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1663859327
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1663859327
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1663859327
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1663859327
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1663859327
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1663859327
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1663859327
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1663859327
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1663859327
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1663859327
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1663859327
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1663859327
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1663859327
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1663859327
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1663859327
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1663859327
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1663859327
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1663859327
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1663859327
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1663859327
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1663859327
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1663859327
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1663859327
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1663859327
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1663859327
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1663859327
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1663859327
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1663859327
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1663859327
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1663859327
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1663859327
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1663859327
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1663859327
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1663859327
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1663859327
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1663859327
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1663859327
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1663859327
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1663859327
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1663859327
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1663859327
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1663859327
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1663859327
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1663859327
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1663859327
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1663859327
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1663859327
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1663859327
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1663859327
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1663859327
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1663859327
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1663859327
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1663859327
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1663859327
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1663859327
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1663859327
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1663859327
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1663859327
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1663859327
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1663859327
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1663859327
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1663859327
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1663859327
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1663859327
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1663859327
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1663859327
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1663859327
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1663859327
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1663859327
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1663859327
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1663859327
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1663859327
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1663859327
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1663859327
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1663859327
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1663859327
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1663859327
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1663859327
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1663859327
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1663859327
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1663859327
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1663859327
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1663859327
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1663859327
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1663859327
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1663859327
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1663859327
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1663859327
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1663859327
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1663859327
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1663859327
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1663859327
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1663859327
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1663859327
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1663859327
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1663859327
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1663859327
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1663859327
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1663859327
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1663859327
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1663859327
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1663859327
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1663859327
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1663859327
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1663859327
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1663859327
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1663859327
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1663859327
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1663859327
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1663859327
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1663859327
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1663859327
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1663859327
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1663859327
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1663859327
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1663859327
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1663859327
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1663859327
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1663859327
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1663859327
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1663859327
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1663859327
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1663859327
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1663859327
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1663859327
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1663859327
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1663859327
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1663859327
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1663859327
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1663859327
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1663859327
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1663859327
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1663859327
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1663859327
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1663859327
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1663859327
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1663859327
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1663859327
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1663859327
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1663859327
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1663859327
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1663859327
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1663859327
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1663859327
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1663859327
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1663859327
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1663859327
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1663859327
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1663859327
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1663859327
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1663859327
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1663859327
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1663859327
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1663859327
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1663859327
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1663859327
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1663859327
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1663859327
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1663859327
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1663859327
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1663859327
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1663859327
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1663859327
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1663859327
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1663859327
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1663859327
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1663859327
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1663859327
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1663859327
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1663859327
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1663859327
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1663859327
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1663859327
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1663859327
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1663859327
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1663859327
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1663859327
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1663859327
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1663859327
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1663859327
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1663859327
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1663859327
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1663859327
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1663859327
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1663859327
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1663859327
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1663859327
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1663859327
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1663859327
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1663859327
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1663859327
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1663859327
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1663859327
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1663859327
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1663859327
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1663859327
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1663859327
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1663859327
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1663859327
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1663859327
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1663859327
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1663859327
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1663859327
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1663859327
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1663859327
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1663859327
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1663859327
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1663859327
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1663859327
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1663859327
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1663859327
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1663859327
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1663859327
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1663859327
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1663859327
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1663859327
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1663859327
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1663859327
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1663859327
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1663859327
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1663859327
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1663859327
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1663859327
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1663859327
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1663859327
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1663859327
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1663859327
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1663859327
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1663859327
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1663859327
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1663859327
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1663859327
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1663859327
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1663859327
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1663859327
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1663859327
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1663859327
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1663859327
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1663859327
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1663859327
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1663859327
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1663859327
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1663859327
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1663859327
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1663859327
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1663859327
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1663859327
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1663859327
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1663859327
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1663859327
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1663859327
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1663859327
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1663859327
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1663859327
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1663859327
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1663859327
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1663859327
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1663859327
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1663859327
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1663859327
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1663859327
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1663859327
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1663859327
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1663859327
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1663859327
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1663859327
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1663859327
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1663859327
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1663859327
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1663859327
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1663859327
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1663859327
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1663859327
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1663859327
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1663859327
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1663859327
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1663859327
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1663859327
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1663859327
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1663859327
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1663859327
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1663859327
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1663859327
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1663859327
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1663859327
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1663859327
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1663859327
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1663859327
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1663859327
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1663859327
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1663859327
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1663859327
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1663859327
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1663859327
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1663859327
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_1 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 2576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_2
timestamp 1663859327
transform -1 0 9968 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_3
timestamp 1663859327
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_4
timestamp 1663859327
transform -1 0 2128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_5
timestamp 1663859327
transform -1 0 2128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_6
timestamp 1663859327
transform 1 0 47824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_7
timestamp 1663859327
transform -1 0 2128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_8
timestamp 1663859327
transform -1 0 2128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_9
timestamp 1663859327
transform 1 0 47824 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_10
timestamp 1663859327
transform 1 0 47824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_11
timestamp 1663859327
transform -1 0 42896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_12
timestamp 1663859327
transform 1 0 47824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_13
timestamp 1663859327
transform -1 0 2128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_14
timestamp 1663859327
transform -1 0 2128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_15
timestamp 1663859327
transform -1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_16
timestamp 1663859327
transform -1 0 2128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_17
timestamp 1663859327
transform -1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_18
timestamp 1663859327
transform -1 0 20720 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_19
timestamp 1663859327
transform -1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_20
timestamp 1663859327
transform -1 0 2128 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_21
timestamp 1663859327
transform -1 0 2128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_22
timestamp 1663859327
transform -1 0 2800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_23
timestamp 1663859327
transform -1 0 43568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_24
timestamp 1663859327
transform -1 0 33488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_25
timestamp 1663859327
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_26
timestamp 1663859327
transform 1 0 47824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_27
timestamp 1663859327
transform -1 0 3248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_28
timestamp 1663859327
transform -1 0 2128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_29
timestamp 1663859327
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_30
timestamp 1663859327
transform -1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_31
timestamp 1663859327
transform -1 0 2128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_32
timestamp 1663859327
transform 1 0 47824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_33
timestamp 1663859327
transform -1 0 29568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_34
timestamp 1663859327
transform -1 0 40208 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_35
timestamp 1663859327
transform -1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_36
timestamp 1663859327
transform -1 0 27440 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_37
timestamp 1663859327
transform -1 0 41328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_38
timestamp 1663859327
transform -1 0 2128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_39
timestamp 1663859327
transform -1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_40
timestamp 1663859327
transform -1 0 2128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_41
timestamp 1663859327
transform 1 0 47824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_42
timestamp 1663859327
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_43
timestamp 1663859327
transform 1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_44
timestamp 1663859327
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_45
timestamp 1663859327
transform -1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_46
timestamp 1663859327
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_47
timestamp 1663859327
transform -1 0 2128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_48
timestamp 1663859327
transform -1 0 2128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_49
timestamp 1663859327
transform 1 0 47824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_50
timestamp 1663859327
transform -1 0 44240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_51
timestamp 1663859327
transform -1 0 2128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_52
timestamp 1663859327
transform 1 0 47824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_53
timestamp 1663859327
transform -1 0 22064 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_54
timestamp 1663859327
transform -1 0 13888 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_55
timestamp 1663859327
transform -1 0 18704 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_56
timestamp 1663859327
transform -1 0 14672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_57
timestamp 1663859327
transform 1 0 47824 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_58
timestamp 1663859327
transform 1 0 47824 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_59
timestamp 1663859327
transform 1 0 47824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_60
timestamp 1663859327
transform -1 0 3920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_61
timestamp 1663859327
transform -1 0 46256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_62
timestamp 1663859327
transform 1 0 47824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_63
timestamp 1663859327
transform -1 0 2128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_64
timestamp 1663859327
transform -1 0 2128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_65
timestamp 1663859327
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_66
timestamp 1663859327
transform 1 0 47824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_67
timestamp 1663859327
transform 1 0 47824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_68
timestamp 1663859327
transform -1 0 2128 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_69
timestamp 1663859327
transform 1 0 47152 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_70
timestamp 1663859327
transform -1 0 2800 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_71
timestamp 1663859327
transform -1 0 7952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_72
timestamp 1663859327
transform -1 0 2128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_73
timestamp 1663859327
transform -1 0 2128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_74
timestamp 1663859327
transform -1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_75
timestamp 1663859327
transform 1 0 47824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_76
timestamp 1663859327
transform -1 0 38192 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal2 s 23520 49200 23632 49800 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 49728 49200 49840 49800 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 24192 200 24304 800 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 11424 49200 11536 49800 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 49056 200 49168 800 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 49200 43008 49800 43120 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 36960 200 37072 800 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 12096 200 12208 800 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 200 47712 800 47824 0 FreeSans 448 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 18816 200 18928 800 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30912 49200 31024 49800 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 200 1344 800 1456 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 33600 200 33712 800 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 200 31584 800 31696 0 FreeSans 448 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal3 s 49200 20160 49800 20272 0 FreeSans 448 0 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 49200 46368 49800 46480 0 FreeSans 448 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 200 4704 800 4816 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 40992 49200 41104 49800 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 200 40320 800 40432 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 49200 14784 49800 14896 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 49200 40992 49800 41104 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 47712 200 47824 800 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 29568 200 29680 800 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 49200 4032 49800 4144 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 14784 49200 14896 49800 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 10080 200 10192 800 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 25536 49200 25648 49800 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 46368 49200 46480 49800 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 200 12096 800 12208 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 16128 49200 16240 49800 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 49200 45024 49800 45136 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 49200 25536 49800 25648 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 28896 49200 29008 49800 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 6720 200 6832 800 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 45024 49200 45136 49800 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 49200 34384 49800 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 6048 49200 6160 49800 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 49200 48384 49800 48496 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 15456 200 15568 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 200 8736 800 8848 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 49200 34272 49800 34384 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 200 34944 800 35056 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 200 18816 800 18928 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 49200 11424 49800 11536 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 43680 200 43792 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal3 s 200 24192 800 24304 0 FreeSans 448 0 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal3 s 49200 26880 49800 26992 0 FreeSans 448 0 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 21504 49200 21616 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 12768 49200 12880 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 26880 49200 26992 49800 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 18144 49200 18256 49800 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 14112 200 14224 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal3 s 49200 12768 49800 12880 0 FreeSans 448 0 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal3 s 49200 6048 49800 6160 0 FreeSans 448 0 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 49200 32256 49800 32368 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 3360 200 3472 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 45696 200 45808 800 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 49200 9408 49800 9520 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 200 29568 800 29680 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 200 3360 800 3472 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 40320 200 40432 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 20832 200 20944 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 49200 16800 49800 16912 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 49200 37632 49800 37744 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 200 38304 800 38416 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 49200 2016 49800 2128 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 200 45696 800 45808 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 7392 49200 7504 49800 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 200 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 200 6720 800 6832 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 4704 200 4816 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 200 20832 800 20944 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 49200 672 49800 784 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 49200 28896 49800 29008 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 49200 18144 49800 18256 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 38304 200 38416 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 200 36960 800 37072 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 200 28224 800 28336 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 200 26208 800 26320 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 49200 21504 49800 21616 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 49200 35616 49800 35728 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 42336 200 42448 800 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal3 s 49200 39648 49800 39760 0 FreeSans 448 0 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 672 49200 784 49800 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal3 s 200 10080 800 10192 0 FreeSans 448 0 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 26208 200 26320 800 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 31584 200 31696 800 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 4032 49200 4144 49800 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 20160 49200 20272 49800 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35616 49200 35728 49800 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal3 s 200 43680 800 43792 0 FreeSans 448 0 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 200 22848 800 22960 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 1344 200 1456 800 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 43008 49200 43120 49800 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 32256 49200 32368 49800 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 22848 200 22960 800 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 48384 49200 48496 49800 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 49200 7392 49800 7504 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 200 49056 800 49168 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 200 17472 800 17584 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 8736 200 8848 800 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 17472 200 17584 800 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 200 15456 800 15568 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 49200 30912 49800 31024 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 28224 200 28336 800 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 39648 49200 39760 49800 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 37632 49200 37744 49800 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 2016 49200 2128 49800 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 9408 49200 9520 49800 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 34944 200 35056 800 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 200 14112 800 14224 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 200 42336 800 42448 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 49200 23520 49800 23632 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vccd1
rlabel metal1 24976 45472 24976 45472 0 vssd1
rlabel metal2 2184 45752 2184 45752 0 net1
rlabel metal2 48104 35952 48104 35952 0 net10
rlabel metal2 42392 2030 42392 2030 0 net11
rlabel metal2 48104 40096 48104 40096 0 net12
rlabel metal2 1848 47320 1848 47320 0 net13
rlabel metal3 1302 10136 1302 10136 0 net14
rlabel metal2 26264 2030 26264 2030 0 net15
rlabel metal2 56 2590 56 2590 0 net16
rlabel metal2 4200 45752 4200 45752 0 net17
rlabel metal2 20328 45752 20328 45752 0 net18
rlabel metal2 35784 45752 35784 45752 0 net19
rlabel metal2 9576 45752 9576 45752 0 net2
rlabel metal3 1302 43736 1302 43736 0 net20
rlabel metal3 1302 22904 1302 22904 0 net21
rlabel metal2 1400 2030 1400 2030 0 net22
rlabel metal2 43176 45752 43176 45752 0 net23
rlabel metal2 33208 46088 33208 46088 0 net24
rlabel metal2 22904 2030 22904 2030 0 net25
rlabel metal2 48272 45752 48272 45752 0 net26
rlabel metal2 2968 46368 2968 46368 0 net27
rlabel metal3 1302 17528 1302 17528 0 net28
rlabel metal2 8792 1246 8792 1246 0 net29
rlabel metal2 35000 2030 35000 2030 0 net3
rlabel metal2 17528 2030 17528 2030 0 net30
rlabel metal3 1302 15512 1302 15512 0 net31
rlabel metal2 48104 31248 48104 31248 0 net32
rlabel metal2 28280 2030 28280 2030 0 net33
rlabel metal2 39816 45752 39816 45752 0 net34
rlabel metal2 15512 2030 15512 2030 0 net35
rlabel metal2 27048 45752 27048 45752 0 net36
rlabel metal2 40376 1302 40376 1302 0 net37
rlabel metal3 1302 6776 1302 6776 0 net38
rlabel metal2 4760 2030 4760 2030 0 net39
rlabel metal3 1302 14168 1302 14168 0 net4
rlabel metal3 1302 20888 1302 20888 0 net40
rlabel metal2 48104 2016 48104 2016 0 net41
rlabel metal2 48104 29232 48104 29232 0 net42
rlabel metal2 48104 18368 48104 18368 0 net43
rlabel metal2 38360 2030 38360 2030 0 net44
rlabel metal3 1302 8792 1302 8792 0 net45
rlabel metal2 48104 34496 48104 34496 0 net46
rlabel metal3 1302 35000 1302 35000 0 net47
rlabel metal3 1302 18872 1302 18872 0 net48
rlabel metal2 48104 11872 48104 11872 0 net49
rlabel metal3 1302 42392 1302 42392 0 net5
rlabel metal2 43736 2030 43736 2030 0 net50
rlabel metal3 1302 24248 1302 24248 0 net51
rlabel metal2 48104 26880 48104 26880 0 net52
rlabel metal2 21672 45752 21672 45752 0 net53
rlabel metal3 13216 45752 13216 45752 0 net54
rlabel metal2 18312 45752 18312 45752 0 net55
rlabel metal2 14168 2030 14168 2030 0 net56
rlabel metal3 48706 12824 48706 12824 0 net57
rlabel metal2 48104 6272 48104 6272 0 net58
rlabel metal2 48104 32480 48104 32480 0 net59
rlabel metal2 48104 23632 48104 23632 0 net6
rlabel metal2 3416 2030 3416 2030 0 net60
rlabel metal2 45752 2030 45752 2030 0 net61
rlabel metal2 48104 9520 48104 9520 0 net62
rlabel metal3 1302 29624 1302 29624 0 net63
rlabel metal2 1848 3360 1848 3360 0 net64
rlabel metal2 20888 1246 20888 1246 0 net65
rlabel metal2 48104 17136 48104 17136 0 net66
rlabel metal2 48104 37744 48104 37744 0 net67
rlabel metal3 1302 38360 1302 38360 0 net68
rlabel metal2 47432 2688 47432 2688 0 net69
rlabel metal3 1302 28280 1302 28280 0 net7
rlabel metal2 2520 45528 2520 45528 0 net70
rlabel metal2 7560 45752 7560 45752 0 net71
rlabel metal3 1302 32984 1302 32984 0 net72
rlabel metal3 1302 37016 1302 37016 0 net73
rlabel metal2 31640 2030 31640 2030 0 net74
rlabel metal2 48104 7728 48104 7728 0 net75
rlabel metal2 37800 45752 37800 45752 0 net76
rlabel metal3 1302 26264 1302 26264 0 net8
rlabel metal2 48104 21840 48104 21840 0 net9
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
